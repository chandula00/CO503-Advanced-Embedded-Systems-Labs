// SoC.v

// Generated using ACDS version 13.1 162 at 2024.05.16.18:42:20

`timescale 1 ps / 1 ps
module SoC (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] mm_interconnect_0_onchip_instruction_memory1_s1_writedata;  // mm_interconnect_0:onchip_instruction_memory1_s1_writedata -> onchip_instruction_memory1:writedata
	wire  [13:0] mm_interconnect_0_onchip_instruction_memory1_s1_address;    // mm_interconnect_0:onchip_instruction_memory1_s1_address -> onchip_instruction_memory1:address
	wire         mm_interconnect_0_onchip_instruction_memory1_s1_chipselect; // mm_interconnect_0:onchip_instruction_memory1_s1_chipselect -> onchip_instruction_memory1:chipselect
	wire         mm_interconnect_0_onchip_instruction_memory1_s1_clken;      // mm_interconnect_0:onchip_instruction_memory1_s1_clken -> onchip_instruction_memory1:clken
	wire         mm_interconnect_0_onchip_instruction_memory1_s1_write;      // mm_interconnect_0:onchip_instruction_memory1_s1_write -> onchip_instruction_memory1:write
	wire  [31:0] mm_interconnect_0_onchip_instruction_memory1_s1_readdata;   // onchip_instruction_memory1:readdata -> mm_interconnect_0:onchip_instruction_memory1_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_instruction_memory1_s1_byteenable; // mm_interconnect_0:onchip_instruction_memory1_s1_byteenable -> onchip_instruction_memory1:byteenable
	wire         cpu0_instruction_master_waitrequest;                        // mm_interconnect_0:cpu0_instruction_master_waitrequest -> cpu0:i_waitrequest
	wire  [18:0] cpu0_instruction_master_address;                            // cpu0:i_address -> mm_interconnect_0:cpu0_instruction_master_address
	wire         cpu0_instruction_master_read;                               // cpu0:i_read -> mm_interconnect_0:cpu0_instruction_master_read
	wire  [31:0] cpu0_instruction_master_readdata;                           // mm_interconnect_0:cpu0_instruction_master_readdata -> cpu0:i_readdata
	wire  [31:0] mm_interconnect_0_onchip_instruction_memory0_s1_writedata;  // mm_interconnect_0:onchip_instruction_memory0_s1_writedata -> onchip_instruction_memory0:writedata
	wire  [13:0] mm_interconnect_0_onchip_instruction_memory0_s1_address;    // mm_interconnect_0:onchip_instruction_memory0_s1_address -> onchip_instruction_memory0:address
	wire         mm_interconnect_0_onchip_instruction_memory0_s1_chipselect; // mm_interconnect_0:onchip_instruction_memory0_s1_chipselect -> onchip_instruction_memory0:chipselect
	wire         mm_interconnect_0_onchip_instruction_memory0_s1_clken;      // mm_interconnect_0:onchip_instruction_memory0_s1_clken -> onchip_instruction_memory0:clken
	wire         mm_interconnect_0_onchip_instruction_memory0_s1_write;      // mm_interconnect_0:onchip_instruction_memory0_s1_write -> onchip_instruction_memory0:write
	wire  [31:0] mm_interconnect_0_onchip_instruction_memory0_s1_readdata;   // onchip_instruction_memory0:readdata -> mm_interconnect_0:onchip_instruction_memory0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_instruction_memory0_s1_byteenable; // mm_interconnect_0:onchip_instruction_memory0_s1_byteenable -> onchip_instruction_memory0:byteenable
	wire         mm_interconnect_0_jtag_uart0_avalon_jtag_slave_waitrequest; // jtag_uart0:av_waitrequest -> mm_interconnect_0:jtag_uart0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart0_avalon_jtag_slave_writedata -> jtag_uart0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart0_avalon_jtag_slave_address -> jtag_uart0:av_address
	wire         mm_interconnect_0_jtag_uart0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart0_avalon_jtag_slave_chipselect -> jtag_uart0:av_chipselect
	wire         mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart0_avalon_jtag_slave_write -> jtag_uart0:av_write_n
	wire         mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart0_avalon_jtag_slave_read -> jtag_uart0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart0_avalon_jtag_slave_readdata;    // jtag_uart0:av_readdata -> mm_interconnect_0:jtag_uart0_avalon_jtag_slave_readdata
	wire         cpu0_data_master_waitrequest;                               // mm_interconnect_0:cpu0_data_master_waitrequest -> cpu0:d_waitrequest
	wire  [31:0] cpu0_data_master_writedata;                                 // cpu0:d_writedata -> mm_interconnect_0:cpu0_data_master_writedata
	wire  [18:0] cpu0_data_master_address;                                   // cpu0:d_address -> mm_interconnect_0:cpu0_data_master_address
	wire         cpu0_data_master_write;                                     // cpu0:d_write -> mm_interconnect_0:cpu0_data_master_write
	wire         cpu0_data_master_read;                                      // cpu0:d_read -> mm_interconnect_0:cpu0_data_master_read
	wire  [31:0] cpu0_data_master_readdata;                                  // mm_interconnect_0:cpu0_data_master_readdata -> cpu0:d_readdata
	wire         cpu0_data_master_debugaccess;                               // cpu0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu0_data_master_debugaccess
	wire   [3:0] cpu0_data_master_byteenable;                                // cpu0:d_byteenable -> mm_interconnect_0:cpu0_data_master_byteenable
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;              // mm_interconnect_0:sysId_control_slave_address -> sysId:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;             // sysId:readdata -> mm_interconnect_0:sysId_control_slave_readdata
	wire  [15:0] mm_interconnect_0_timer0_s1_writedata;                      // mm_interconnect_0:timer0_s1_writedata -> timer0:writedata
	wire   [2:0] mm_interconnect_0_timer0_s1_address;                        // mm_interconnect_0:timer0_s1_address -> timer0:address
	wire         mm_interconnect_0_timer0_s1_chipselect;                     // mm_interconnect_0:timer0_s1_chipselect -> timer0:chipselect
	wire         mm_interconnect_0_timer0_s1_write;                          // mm_interconnect_0:timer0_s1_write -> timer0:write_n
	wire  [15:0] mm_interconnect_0_timer0_s1_readdata;                       // timer0:readdata -> mm_interconnect_0:timer0_s1_readdata
	wire         mm_interconnect_0_cpu0_jtag_debug_module_waitrequest;       // cpu0:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu0_jtag_debug_module_writedata;         // mm_interconnect_0:cpu0_jtag_debug_module_writedata -> cpu0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu0_jtag_debug_module_address;           // mm_interconnect_0:cpu0_jtag_debug_module_address -> cpu0:jtag_debug_module_address
	wire         mm_interconnect_0_cpu0_jtag_debug_module_write;             // mm_interconnect_0:cpu0_jtag_debug_module_write -> cpu0:jtag_debug_module_write
	wire         mm_interconnect_0_cpu0_jtag_debug_module_read;              // mm_interconnect_0:cpu0_jtag_debug_module_read -> cpu0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu0_jtag_debug_module_readdata;          // cpu0:jtag_debug_module_readdata -> mm_interconnect_0:cpu0_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu0_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu0_jtag_debug_module_debugaccess -> cpu0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu0_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu0_jtag_debug_module_byteenable -> cpu0:jtag_debug_module_byteenable
	wire         cpu1_instruction_master_waitrequest;                        // mm_interconnect_0:cpu1_instruction_master_waitrequest -> cpu1:i_waitrequest
	wire  [18:0] cpu1_instruction_master_address;                            // cpu1:i_address -> mm_interconnect_0:cpu1_instruction_master_address
	wire         cpu1_instruction_master_read;                               // cpu1:i_read -> mm_interconnect_0:cpu1_instruction_master_read
	wire  [31:0] cpu1_instruction_master_readdata;                           // mm_interconnect_0:cpu1_instruction_master_readdata -> cpu1:i_readdata
	wire  [15:0] mm_interconnect_0_timer1_s1_writedata;                      // mm_interconnect_0:timer1_s1_writedata -> timer1:writedata
	wire   [2:0] mm_interconnect_0_timer1_s1_address;                        // mm_interconnect_0:timer1_s1_address -> timer1:address
	wire         mm_interconnect_0_timer1_s1_chipselect;                     // mm_interconnect_0:timer1_s1_chipselect -> timer1:chipselect
	wire         mm_interconnect_0_timer1_s1_write;                          // mm_interconnect_0:timer1_s1_write -> timer1:write_n
	wire  [15:0] mm_interconnect_0_timer1_s1_readdata;                       // timer1:readdata -> mm_interconnect_0:timer1_s1_readdata
	wire         mm_interconnect_0_fifo_mem_out_waitrequest;                 // fifo_mem:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_mem_out_waitrequest
	wire         mm_interconnect_0_fifo_mem_out_read;                        // mm_interconnect_0:fifo_mem_out_read -> fifo_mem:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_mem_out_readdata;                    // fifo_mem:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_mem_out_readdata
	wire         mm_interconnect_0_fifo_mem_in_waitrequest;                  // fifo_mem:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_mem_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_mem_in_writedata;                    // mm_interconnect_0:fifo_mem_in_writedata -> fifo_mem:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_mem_in_write;                        // mm_interconnect_0:fifo_mem_in_write -> fifo_mem:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo_mem_in_csr_writedata;                // mm_interconnect_0:fifo_mem_in_csr_writedata -> fifo_mem:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_mem_in_csr_address;                  // mm_interconnect_0:fifo_mem_in_csr_address -> fifo_mem:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_mem_in_csr_write;                    // mm_interconnect_0:fifo_mem_in_csr_write -> fifo_mem:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_mem_in_csr_read;                     // mm_interconnect_0:fifo_mem_in_csr_read -> fifo_mem:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_mem_in_csr_readdata;                 // fifo_mem:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_mem_in_csr_readdata
	wire         mm_interconnect_0_cpu1_jtag_debug_module_waitrequest;       // cpu1:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu1_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu1_jtag_debug_module_writedata;         // mm_interconnect_0:cpu1_jtag_debug_module_writedata -> cpu1:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu1_jtag_debug_module_address;           // mm_interconnect_0:cpu1_jtag_debug_module_address -> cpu1:jtag_debug_module_address
	wire         mm_interconnect_0_cpu1_jtag_debug_module_write;             // mm_interconnect_0:cpu1_jtag_debug_module_write -> cpu1:jtag_debug_module_write
	wire         mm_interconnect_0_cpu1_jtag_debug_module_read;              // mm_interconnect_0:cpu1_jtag_debug_module_read -> cpu1:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu1_jtag_debug_module_readdata;          // cpu1:jtag_debug_module_readdata -> mm_interconnect_0:cpu1_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu1_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu1_jtag_debug_module_debugaccess -> cpu1:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu1_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu1_jtag_debug_module_byteenable -> cpu1:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_data_memory_cpu1_s1_writedata;     // mm_interconnect_0:onchip_data_memory_cpu1_s1_writedata -> onchip_data_memory_cpu1:writedata
	wire  [14:0] mm_interconnect_0_onchip_data_memory_cpu1_s1_address;       // mm_interconnect_0:onchip_data_memory_cpu1_s1_address -> onchip_data_memory_cpu1:address
	wire         mm_interconnect_0_onchip_data_memory_cpu1_s1_chipselect;    // mm_interconnect_0:onchip_data_memory_cpu1_s1_chipselect -> onchip_data_memory_cpu1:chipselect
	wire         mm_interconnect_0_onchip_data_memory_cpu1_s1_clken;         // mm_interconnect_0:onchip_data_memory_cpu1_s1_clken -> onchip_data_memory_cpu1:clken
	wire         mm_interconnect_0_onchip_data_memory_cpu1_s1_write;         // mm_interconnect_0:onchip_data_memory_cpu1_s1_write -> onchip_data_memory_cpu1:write
	wire  [31:0] mm_interconnect_0_onchip_data_memory_cpu1_s1_readdata;      // onchip_data_memory_cpu1:readdata -> mm_interconnect_0:onchip_data_memory_cpu1_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_data_memory_cpu1_s1_byteenable;    // mm_interconnect_0:onchip_data_memory_cpu1_s1_byteenable -> onchip_data_memory_cpu1:byteenable
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest; // jtag_uart1:av_waitrequest -> mm_interconnect_0:jtag_uart1_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_writedata -> jtag_uart1:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_address -> jtag_uart1:av_address
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_chipselect -> jtag_uart1:av_chipselect
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_write -> jtag_uart1:av_write_n
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_read -> jtag_uart1:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata;    // jtag_uart1:av_readdata -> mm_interconnect_0:jtag_uart1_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_onchip_data_memory_cpu0_s1_writedata;     // mm_interconnect_0:onchip_data_memory_cpu0_s1_writedata -> onchip_data_memory_cpu0:writedata
	wire  [14:0] mm_interconnect_0_onchip_data_memory_cpu0_s1_address;       // mm_interconnect_0:onchip_data_memory_cpu0_s1_address -> onchip_data_memory_cpu0:address
	wire         mm_interconnect_0_onchip_data_memory_cpu0_s1_chipselect;    // mm_interconnect_0:onchip_data_memory_cpu0_s1_chipselect -> onchip_data_memory_cpu0:chipselect
	wire         mm_interconnect_0_onchip_data_memory_cpu0_s1_clken;         // mm_interconnect_0:onchip_data_memory_cpu0_s1_clken -> onchip_data_memory_cpu0:clken
	wire         mm_interconnect_0_onchip_data_memory_cpu0_s1_write;         // mm_interconnect_0:onchip_data_memory_cpu0_s1_write -> onchip_data_memory_cpu0:write
	wire  [31:0] mm_interconnect_0_onchip_data_memory_cpu0_s1_readdata;      // onchip_data_memory_cpu0:readdata -> mm_interconnect_0:onchip_data_memory_cpu0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_data_memory_cpu0_s1_byteenable;    // mm_interconnect_0:onchip_data_memory_cpu0_s1_byteenable -> onchip_data_memory_cpu0:byteenable
	wire         cpu1_data_master_waitrequest;                               // mm_interconnect_0:cpu1_data_master_waitrequest -> cpu1:d_waitrequest
	wire  [31:0] cpu1_data_master_writedata;                                 // cpu1:d_writedata -> mm_interconnect_0:cpu1_data_master_writedata
	wire  [18:0] cpu1_data_master_address;                                   // cpu1:d_address -> mm_interconnect_0:cpu1_data_master_address
	wire         cpu1_data_master_write;                                     // cpu1:d_write -> mm_interconnect_0:cpu1_data_master_write
	wire         cpu1_data_master_read;                                      // cpu1:d_read -> mm_interconnect_0:cpu1_data_master_read
	wire  [31:0] cpu1_data_master_readdata;                                  // mm_interconnect_0:cpu1_data_master_readdata -> cpu1:d_readdata
	wire         cpu1_data_master_debugaccess;                               // cpu1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu1_data_master_debugaccess
	wire   [3:0] cpu1_data_master_byteenable;                                // cpu1:d_byteenable -> mm_interconnect_0:cpu1_data_master_byteenable
	wire         irq_mapper_receiver0_irq;                                   // timer0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // jtag_uart0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu0_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu0:d_irq
	wire         irq_mapper_001_receiver0_irq;                               // timer1:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                               // jtag_uart1:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu1_d_irq_irq;                                             // irq_mapper_001:sender_irq -> cpu1:d_irq
	wire         irq_mapper_receiver2_irq;                                   // fifo_mem:wrclk_control_slave_irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq]
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [cpu0:reset_n, irq_mapper:reset, jtag_uart0:rst_n, mm_interconnect_0:cpu0_reset_n_reset_bridge_in_reset_reset, onchip_data_memory_cpu0:reset, onchip_instruction_memory0:reset, rst_translator:in_reset, timer0:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [cpu0:reset_req, onchip_data_memory_cpu0:reset_req, onchip_instruction_memory0:reset_req, rst_translator:reset_req_in]
	wire         cpu0_jtag_debug_module_reset_reset;                         // cpu0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [cpu1:reset_n, irq_mapper_001:reset, jtag_uart1:rst_n, mm_interconnect_0:cpu1_reset_n_reset_bridge_in_reset_reset, onchip_data_memory_cpu1:reset, onchip_instruction_memory1:reset, rst_translator_001:in_reset, timer1:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> [cpu1:reset_req, onchip_data_memory_cpu1:reset_req, onchip_instruction_memory1:reset_req, rst_translator_001:reset_req_in]
	wire         cpu1_jtag_debug_module_reset_reset;                         // cpu1:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_002:reset_in2]
	wire         rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [fifo_mem:reset_n, mm_interconnect_0:sysId_reset_reset_bridge_in_reset_reset, sysId:reset_n]

	SoC_cpu0 cpu0 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (cpu0_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu0_data_master_read),                                //                          .read
		.d_readdata                            (cpu0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu0_data_master_write),                               //                          .write
		.d_writedata                           (cpu0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu0_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	SoC_cpu1 cpu1 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                  //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),               //                          .reset_req
		.d_address                             (cpu1_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu1_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu1_data_master_read),                                //                          .read
		.d_readdata                            (cpu1_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu1_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu1_data_master_write),                               //                          .write
		.d_writedata                           (cpu1_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu1_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu1_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu1_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu1_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu1_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu1_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu1_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu1_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu1_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu1_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu1_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu1_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu1_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu1_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu1_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	SoC_timer0 timer0 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                //   irq.irq
	);

	SoC_timer0 timer1 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    // reset.reset_n
		.address    (mm_interconnect_0_timer1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)            //   irq.irq
	);

	SoC_jtag_uart0 jtag_uart0 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                            //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                    //               irq.irq
	);

	SoC_jtag_uart0 jtag_uart1 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                //               irq.irq
	);

	SoC_onchip_instruction_memory0 onchip_instruction_memory0 (
		.clk        (clk_clk),                                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_instruction_memory0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_instruction_memory0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_instruction_memory0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_instruction_memory0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_instruction_memory0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_instruction_memory0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_instruction_memory0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                          //       .reset_req
	);

	SoC_onchip_instruction_memory1 onchip_instruction_memory1 (
		.clk        (clk_clk),                                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_instruction_memory1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_instruction_memory1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_instruction_memory1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_instruction_memory1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_instruction_memory1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_instruction_memory1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_instruction_memory1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                         // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)                      //       .reset_req
	);

	SoC_onchip_data_memory_cpu0 onchip_data_memory_cpu0 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (mm_interconnect_0_onchip_data_memory_cpu0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_data_memory_cpu0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_data_memory_cpu0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_data_memory_cpu0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_data_memory_cpu0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_data_memory_cpu0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_data_memory_cpu0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                       //       .reset_req
	);

	SoC_sysId sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	SoC_fifo_mem fifo_mem (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_002_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_mem_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_mem_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_mem_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_mem_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_mem_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_mem_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_mem_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_mem_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_mem_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_mem_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_mem_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver2_irq)                     //   in_irq.irq
	);

	SoC_onchip_data_memory_cpu1 onchip_data_memory_cpu1 (
		.clk        (clk_clk),                                                 //   clk1.clk
		.address    (mm_interconnect_0_onchip_data_memory_cpu1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_data_memory_cpu1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_data_memory_cpu1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_data_memory_cpu1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_data_memory_cpu1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_data_memory_cpu1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_data_memory_cpu1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                      // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)                   //       .reset_req
	);

	SoC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                            (clk_clk),                                                    //                          clock_clk.clk
		.cpu0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // cpu0_reset_n_reset_bridge_in_reset.reset
		.cpu1_reset_n_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // cpu1_reset_n_reset_bridge_in_reset.reset
		.sysId_reset_reset_bridge_in_reset_reset  (rst_controller_002_reset_out_reset),                         //  sysId_reset_reset_bridge_in_reset.reset
		.cpu0_data_master_address                 (cpu0_data_master_address),                                   //                   cpu0_data_master.address
		.cpu0_data_master_waitrequest             (cpu0_data_master_waitrequest),                               //                                   .waitrequest
		.cpu0_data_master_byteenable              (cpu0_data_master_byteenable),                                //                                   .byteenable
		.cpu0_data_master_read                    (cpu0_data_master_read),                                      //                                   .read
		.cpu0_data_master_readdata                (cpu0_data_master_readdata),                                  //                                   .readdata
		.cpu0_data_master_write                   (cpu0_data_master_write),                                     //                                   .write
		.cpu0_data_master_writedata               (cpu0_data_master_writedata),                                 //                                   .writedata
		.cpu0_data_master_debugaccess             (cpu0_data_master_debugaccess),                               //                                   .debugaccess
		.cpu0_instruction_master_address          (cpu0_instruction_master_address),                            //            cpu0_instruction_master.address
		.cpu0_instruction_master_waitrequest      (cpu0_instruction_master_waitrequest),                        //                                   .waitrequest
		.cpu0_instruction_master_read             (cpu0_instruction_master_read),                               //                                   .read
		.cpu0_instruction_master_readdata         (cpu0_instruction_master_readdata),                           //                                   .readdata
		.cpu1_data_master_address                 (cpu1_data_master_address),                                   //                   cpu1_data_master.address
		.cpu1_data_master_waitrequest             (cpu1_data_master_waitrequest),                               //                                   .waitrequest
		.cpu1_data_master_byteenable              (cpu1_data_master_byteenable),                                //                                   .byteenable
		.cpu1_data_master_read                    (cpu1_data_master_read),                                      //                                   .read
		.cpu1_data_master_readdata                (cpu1_data_master_readdata),                                  //                                   .readdata
		.cpu1_data_master_write                   (cpu1_data_master_write),                                     //                                   .write
		.cpu1_data_master_writedata               (cpu1_data_master_writedata),                                 //                                   .writedata
		.cpu1_data_master_debugaccess             (cpu1_data_master_debugaccess),                               //                                   .debugaccess
		.cpu1_instruction_master_address          (cpu1_instruction_master_address),                            //            cpu1_instruction_master.address
		.cpu1_instruction_master_waitrequest      (cpu1_instruction_master_waitrequest),                        //                                   .waitrequest
		.cpu1_instruction_master_read             (cpu1_instruction_master_read),                               //                                   .read
		.cpu1_instruction_master_readdata         (cpu1_instruction_master_readdata),                           //                                   .readdata
		.cpu0_jtag_debug_module_address           (mm_interconnect_0_cpu0_jtag_debug_module_address),           //             cpu0_jtag_debug_module.address
		.cpu0_jtag_debug_module_write             (mm_interconnect_0_cpu0_jtag_debug_module_write),             //                                   .write
		.cpu0_jtag_debug_module_read              (mm_interconnect_0_cpu0_jtag_debug_module_read),              //                                   .read
		.cpu0_jtag_debug_module_readdata          (mm_interconnect_0_cpu0_jtag_debug_module_readdata),          //                                   .readdata
		.cpu0_jtag_debug_module_writedata         (mm_interconnect_0_cpu0_jtag_debug_module_writedata),         //                                   .writedata
		.cpu0_jtag_debug_module_byteenable        (mm_interconnect_0_cpu0_jtag_debug_module_byteenable),        //                                   .byteenable
		.cpu0_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu0_jtag_debug_module_waitrequest),       //                                   .waitrequest
		.cpu0_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu0_jtag_debug_module_debugaccess),       //                                   .debugaccess
		.cpu1_jtag_debug_module_address           (mm_interconnect_0_cpu1_jtag_debug_module_address),           //             cpu1_jtag_debug_module.address
		.cpu1_jtag_debug_module_write             (mm_interconnect_0_cpu1_jtag_debug_module_write),             //                                   .write
		.cpu1_jtag_debug_module_read              (mm_interconnect_0_cpu1_jtag_debug_module_read),              //                                   .read
		.cpu1_jtag_debug_module_readdata          (mm_interconnect_0_cpu1_jtag_debug_module_readdata),          //                                   .readdata
		.cpu1_jtag_debug_module_writedata         (mm_interconnect_0_cpu1_jtag_debug_module_writedata),         //                                   .writedata
		.cpu1_jtag_debug_module_byteenable        (mm_interconnect_0_cpu1_jtag_debug_module_byteenable),        //                                   .byteenable
		.cpu1_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu1_jtag_debug_module_waitrequest),       //                                   .waitrequest
		.cpu1_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu1_jtag_debug_module_debugaccess),       //                                   .debugaccess
		.fifo_mem_in_write                        (mm_interconnect_0_fifo_mem_in_write),                        //                        fifo_mem_in.write
		.fifo_mem_in_writedata                    (mm_interconnect_0_fifo_mem_in_writedata),                    //                                   .writedata
		.fifo_mem_in_waitrequest                  (mm_interconnect_0_fifo_mem_in_waitrequest),                  //                                   .waitrequest
		.fifo_mem_in_csr_address                  (mm_interconnect_0_fifo_mem_in_csr_address),                  //                    fifo_mem_in_csr.address
		.fifo_mem_in_csr_write                    (mm_interconnect_0_fifo_mem_in_csr_write),                    //                                   .write
		.fifo_mem_in_csr_read                     (mm_interconnect_0_fifo_mem_in_csr_read),                     //                                   .read
		.fifo_mem_in_csr_readdata                 (mm_interconnect_0_fifo_mem_in_csr_readdata),                 //                                   .readdata
		.fifo_mem_in_csr_writedata                (mm_interconnect_0_fifo_mem_in_csr_writedata),                //                                   .writedata
		.fifo_mem_out_read                        (mm_interconnect_0_fifo_mem_out_read),                        //                       fifo_mem_out.read
		.fifo_mem_out_readdata                    (mm_interconnect_0_fifo_mem_out_readdata),                    //                                   .readdata
		.fifo_mem_out_waitrequest                 (mm_interconnect_0_fifo_mem_out_waitrequest),                 //                                   .waitrequest
		.jtag_uart0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_address),     //       jtag_uart0_avalon_jtag_slave.address
		.jtag_uart0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_write),       //                                   .write
		.jtag_uart0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_read),        //                                   .read
		.jtag_uart0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_uart0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_uart0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_uart0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart0_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.jtag_uart1_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address),     //       jtag_uart1_avalon_jtag_slave.address
		.jtag_uart1_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write),       //                                   .write
		.jtag_uart1_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read),        //                                   .read
		.jtag_uart1_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_uart1_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_uart1_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_uart1_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.onchip_data_memory_cpu0_s1_address       (mm_interconnect_0_onchip_data_memory_cpu0_s1_address),       //         onchip_data_memory_cpu0_s1.address
		.onchip_data_memory_cpu0_s1_write         (mm_interconnect_0_onchip_data_memory_cpu0_s1_write),         //                                   .write
		.onchip_data_memory_cpu0_s1_readdata      (mm_interconnect_0_onchip_data_memory_cpu0_s1_readdata),      //                                   .readdata
		.onchip_data_memory_cpu0_s1_writedata     (mm_interconnect_0_onchip_data_memory_cpu0_s1_writedata),     //                                   .writedata
		.onchip_data_memory_cpu0_s1_byteenable    (mm_interconnect_0_onchip_data_memory_cpu0_s1_byteenable),    //                                   .byteenable
		.onchip_data_memory_cpu0_s1_chipselect    (mm_interconnect_0_onchip_data_memory_cpu0_s1_chipselect),    //                                   .chipselect
		.onchip_data_memory_cpu0_s1_clken         (mm_interconnect_0_onchip_data_memory_cpu0_s1_clken),         //                                   .clken
		.onchip_data_memory_cpu1_s1_address       (mm_interconnect_0_onchip_data_memory_cpu1_s1_address),       //         onchip_data_memory_cpu1_s1.address
		.onchip_data_memory_cpu1_s1_write         (mm_interconnect_0_onchip_data_memory_cpu1_s1_write),         //                                   .write
		.onchip_data_memory_cpu1_s1_readdata      (mm_interconnect_0_onchip_data_memory_cpu1_s1_readdata),      //                                   .readdata
		.onchip_data_memory_cpu1_s1_writedata     (mm_interconnect_0_onchip_data_memory_cpu1_s1_writedata),     //                                   .writedata
		.onchip_data_memory_cpu1_s1_byteenable    (mm_interconnect_0_onchip_data_memory_cpu1_s1_byteenable),    //                                   .byteenable
		.onchip_data_memory_cpu1_s1_chipselect    (mm_interconnect_0_onchip_data_memory_cpu1_s1_chipselect),    //                                   .chipselect
		.onchip_data_memory_cpu1_s1_clken         (mm_interconnect_0_onchip_data_memory_cpu1_s1_clken),         //                                   .clken
		.onchip_instruction_memory0_s1_address    (mm_interconnect_0_onchip_instruction_memory0_s1_address),    //      onchip_instruction_memory0_s1.address
		.onchip_instruction_memory0_s1_write      (mm_interconnect_0_onchip_instruction_memory0_s1_write),      //                                   .write
		.onchip_instruction_memory0_s1_readdata   (mm_interconnect_0_onchip_instruction_memory0_s1_readdata),   //                                   .readdata
		.onchip_instruction_memory0_s1_writedata  (mm_interconnect_0_onchip_instruction_memory0_s1_writedata),  //                                   .writedata
		.onchip_instruction_memory0_s1_byteenable (mm_interconnect_0_onchip_instruction_memory0_s1_byteenable), //                                   .byteenable
		.onchip_instruction_memory0_s1_chipselect (mm_interconnect_0_onchip_instruction_memory0_s1_chipselect), //                                   .chipselect
		.onchip_instruction_memory0_s1_clken      (mm_interconnect_0_onchip_instruction_memory0_s1_clken),      //                                   .clken
		.onchip_instruction_memory1_s1_address    (mm_interconnect_0_onchip_instruction_memory1_s1_address),    //      onchip_instruction_memory1_s1.address
		.onchip_instruction_memory1_s1_write      (mm_interconnect_0_onchip_instruction_memory1_s1_write),      //                                   .write
		.onchip_instruction_memory1_s1_readdata   (mm_interconnect_0_onchip_instruction_memory1_s1_readdata),   //                                   .readdata
		.onchip_instruction_memory1_s1_writedata  (mm_interconnect_0_onchip_instruction_memory1_s1_writedata),  //                                   .writedata
		.onchip_instruction_memory1_s1_byteenable (mm_interconnect_0_onchip_instruction_memory1_s1_byteenable), //                                   .byteenable
		.onchip_instruction_memory1_s1_chipselect (mm_interconnect_0_onchip_instruction_memory1_s1_chipselect), //                                   .chipselect
		.onchip_instruction_memory1_s1_clken      (mm_interconnect_0_onchip_instruction_memory1_s1_clken),      //                                   .clken
		.sysId_control_slave_address              (mm_interconnect_0_sysid_control_slave_address),              //                sysId_control_slave.address
		.sysId_control_slave_readdata             (mm_interconnect_0_sysid_control_slave_readdata),             //                                   .readdata
		.timer0_s1_address                        (mm_interconnect_0_timer0_s1_address),                        //                          timer0_s1.address
		.timer0_s1_write                          (mm_interconnect_0_timer0_s1_write),                          //                                   .write
		.timer0_s1_readdata                       (mm_interconnect_0_timer0_s1_readdata),                       //                                   .readdata
		.timer0_s1_writedata                      (mm_interconnect_0_timer0_s1_writedata),                      //                                   .writedata
		.timer0_s1_chipselect                     (mm_interconnect_0_timer0_s1_chipselect),                     //                                   .chipselect
		.timer1_s1_address                        (mm_interconnect_0_timer1_s1_address),                        //                          timer1_s1.address
		.timer1_s1_write                          (mm_interconnect_0_timer1_s1_write),                          //                                   .write
		.timer1_s1_readdata                       (mm_interconnect_0_timer1_s1_readdata),                       //                                   .readdata
		.timer1_s1_writedata                      (mm_interconnect_0_timer1_s1_writedata),                      //                                   .writedata
		.timer1_s1_chipselect                     (mm_interconnect_0_timer1_s1_chipselect)                      //                                   .chipselect
	);

	SoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu0_d_irq_irq)                  //    sender.irq
	);

	SoC_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (cpu1_d_irq_irq)                      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu1_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
