// MSoC.v

// Generated using ACDS version 13.1 162 at 2024.05.29.23:52:55

`timescale 1 ps / 1 ps
module MSoC (
		input  wire        clk_clk,                     //                   clk.clk
		input  wire        reset_reset_n,               //                 reset.reset_n
		output wire [12:0] sdram_controller_wire_addr,  // sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,    //                      .ba
		output wire        sdram_controller_wire_cas_n, //                      .cas_n
		output wire        sdram_controller_wire_cke,   //                      .cke
		output wire        sdram_controller_wire_cs_n,  //                      .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,    //                      .dq
		output wire [3:0]  sdram_controller_wire_dqm,   //                      .dqm
		output wire        sdram_controller_wire_ras_n, //                      .ras_n
		output wire        sdram_controller_wire_we_n,  //                      .we_n
		output wire        pll_c0_clk                   //                pll_c0.clk
	);

	wire         mm_interconnect_0_fifo3to4_out_waitrequest;                 // fifo3to4:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo3to4_out_waitrequest
	wire         mm_interconnect_0_fifo3to4_out_read;                        // mm_interconnect_0:fifo3to4_out_read -> fifo3to4:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo3to4_out_readdata;                    // fifo3to4:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo3to4_out_readdata
	wire         cpu2_data_master_waitrequest;                               // mm_interconnect_0:cpu2_data_master_waitrequest -> cpu2:d_waitrequest
	wire  [31:0] cpu2_data_master_writedata;                                 // cpu2:d_writedata -> mm_interconnect_0:cpu2_data_master_writedata
	wire  [28:0] cpu2_data_master_address;                                   // cpu2:d_address -> mm_interconnect_0:cpu2_data_master_address
	wire         cpu2_data_master_write;                                     // cpu2:d_write -> mm_interconnect_0:cpu2_data_master_write
	wire         cpu2_data_master_read;                                      // cpu2:d_read -> mm_interconnect_0:cpu2_data_master_read
	wire  [31:0] cpu2_data_master_readdata;                                  // mm_interconnect_0:cpu2_data_master_readdata -> cpu2:d_readdata
	wire         cpu2_data_master_debugaccess;                               // cpu2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu2_data_master_debugaccess
	wire   [3:0] cpu2_data_master_byteenable;                                // cpu2:d_byteenable -> mm_interconnect_0:cpu2_data_master_byteenable
	wire         cpu4_instruction_master_waitrequest;                        // mm_interconnect_0:cpu4_instruction_master_waitrequest -> cpu4:i_waitrequest
	wire  [17:0] cpu4_instruction_master_address;                            // cpu4:i_address -> mm_interconnect_0:cpu4_instruction_master_address
	wire         cpu4_instruction_master_read;                               // cpu4:i_read -> mm_interconnect_0:cpu4_instruction_master_read
	wire  [31:0] cpu4_instruction_master_readdata;                           // mm_interconnect_0:cpu4_instruction_master_readdata -> cpu4:i_readdata
	wire  [15:0] mm_interconnect_0_timer4_s1_writedata;                      // mm_interconnect_0:timer4_s1_writedata -> timer4:writedata
	wire   [2:0] mm_interconnect_0_timer4_s1_address;                        // mm_interconnect_0:timer4_s1_address -> timer4:address
	wire         mm_interconnect_0_timer4_s1_chipselect;                     // mm_interconnect_0:timer4_s1_chipselect -> timer4:chipselect
	wire         mm_interconnect_0_timer4_s1_write;                          // mm_interconnect_0:timer4_s1_write -> timer4:write_n
	wire  [15:0] mm_interconnect_0_timer4_s1_readdata;                       // timer4:readdata -> mm_interconnect_0:timer4_s1_readdata
	wire         mm_interconnect_0_fifo1to5_in_waitrequest;                  // fifo1to5:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo1to5_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo1to5_in_writedata;                    // mm_interconnect_0:fifo1to5_in_writedata -> fifo1to5:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo1to5_in_write;                        // mm_interconnect_0:fifo1to5_in_write -> fifo1to5:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo5to6_out_waitrequest;                 // fifo5to6:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo5to6_out_waitrequest
	wire         mm_interconnect_0_fifo5to6_out_read;                        // mm_interconnect_0:fifo5to6_out_read -> fifo5to6:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo5to6_out_readdata;                    // fifo5to6:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo5to6_out_readdata
	wire         mm_interconnect_0_fifo1to4_in_waitrequest;                  // fifo1to4:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo1to4_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo1to4_in_writedata;                    // mm_interconnect_0:fifo1to4_in_writedata -> fifo1to4:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo1to4_in_write;                        // mm_interconnect_0:fifo1to4_in_write -> fifo1to4:avalonmm_write_slave_write
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;          // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;            // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;              // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;           // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire         mm_interconnect_0_sdram_controller_s1_write;                // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire         mm_interconnect_0_sdram_controller_s1_read;                 // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;             // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;        // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;           // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                  // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                    // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_write;                      // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire         mm_interconnect_0_pll_pll_slave_read;                       // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                   // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire         mm_interconnect_0_fifo1to6_out_waitrequest;                 // fifo1to6:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1to6_out_waitrequest
	wire         mm_interconnect_0_fifo1to6_out_read;                        // mm_interconnect_0:fifo1to6_out_read -> fifo1to6:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to6_out_readdata;                    // fifo1to6:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1to6_out_readdata
	wire  [31:0] mm_interconnect_0_mem2_s1_writedata;                        // mm_interconnect_0:mem2_s1_writedata -> mem2:writedata
	wire  [14:0] mm_interconnect_0_mem2_s1_address;                          // mm_interconnect_0:mem2_s1_address -> mem2:address
	wire         mm_interconnect_0_mem2_s1_chipselect;                       // mm_interconnect_0:mem2_s1_chipselect -> mem2:chipselect
	wire         mm_interconnect_0_mem2_s1_clken;                            // mm_interconnect_0:mem2_s1_clken -> mem2:clken
	wire         mm_interconnect_0_mem2_s1_write;                            // mm_interconnect_0:mem2_s1_write -> mem2:write
	wire  [31:0] mm_interconnect_0_mem2_s1_readdata;                         // mem2:readdata -> mm_interconnect_0:mem2_s1_readdata
	wire   [3:0] mm_interconnect_0_mem2_s1_byteenable;                       // mm_interconnect_0:mem2_s1_byteenable -> mem2:byteenable
	wire  [31:0] mm_interconnect_0_fifo1to2a_in_csr_writedata;               // mm_interconnect_0:fifo1to2A_in_csr_writedata -> fifo1to2A:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo1to2a_in_csr_address;                 // mm_interconnect_0:fifo1to2A_in_csr_address -> fifo1to2A:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo1to2a_in_csr_write;                   // mm_interconnect_0:fifo1to2A_in_csr_write -> fifo1to2A:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo1to2a_in_csr_read;                    // mm_interconnect_0:fifo1to2A_in_csr_read -> fifo1to2A:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to2a_in_csr_readdata;                // fifo1to2A:wrclk_control_slave_readdata -> mm_interconnect_0:fifo1to2A_in_csr_readdata
	wire  [15:0] mm_interconnect_0_timer2_s1_writedata;                      // mm_interconnect_0:timer2_s1_writedata -> timer2:writedata
	wire   [2:0] mm_interconnect_0_timer2_s1_address;                        // mm_interconnect_0:timer2_s1_address -> timer2:address
	wire         mm_interconnect_0_timer2_s1_chipselect;                     // mm_interconnect_0:timer2_s1_chipselect -> timer2:chipselect
	wire         mm_interconnect_0_timer2_s1_write;                          // mm_interconnect_0:timer2_s1_write -> timer2:write_n
	wire  [15:0] mm_interconnect_0_timer2_s1_readdata;                       // timer2:readdata -> mm_interconnect_0:timer2_s1_readdata
	wire         mm_interconnect_0_fifo1to5_out_waitrequest;                 // fifo1to5:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1to5_out_waitrequest
	wire         mm_interconnect_0_fifo1to5_out_read;                        // mm_interconnect_0:fifo1to5_out_read -> fifo1to5:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to5_out_readdata;                    // fifo1to5:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1to5_out_readdata
	wire         mm_interconnect_0_fifo4to5_in_waitrequest;                  // fifo4to5:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo4to5_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo4to5_in_writedata;                    // mm_interconnect_0:fifo4to5_in_writedata -> fifo4to5:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo4to5_in_write;                        // mm_interconnect_0:fifo4to5_in_write -> fifo4to5:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo1to2c_out_waitrequest;                // fifo1to2C:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1to2C_out_waitrequest
	wire         mm_interconnect_0_fifo1to2c_out_read;                       // mm_interconnect_0:fifo1to2C_out_read -> fifo1to2C:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to2c_out_readdata;                   // fifo1to2C:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1to2C_out_readdata
	wire         mm_interconnect_0_fifo3to4_in_waitrequest;                  // fifo3to4:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo3to4_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo3to4_in_writedata;                    // mm_interconnect_0:fifo3to4_in_writedata -> fifo3to4:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo3to4_in_write;                        // mm_interconnect_0:fifo3to4_in_write -> fifo3to4:avalonmm_write_slave_write
	wire         cpu1_data_master_waitrequest;                               // mm_interconnect_0:cpu1_data_master_waitrequest -> cpu1:d_waitrequest
	wire  [31:0] cpu1_data_master_writedata;                                 // cpu1:d_writedata -> mm_interconnect_0:cpu1_data_master_writedata
	wire  [28:0] cpu1_data_master_address;                                   // cpu1:d_address -> mm_interconnect_0:cpu1_data_master_address
	wire         cpu1_data_master_write;                                     // cpu1:d_write -> mm_interconnect_0:cpu1_data_master_write
	wire         cpu1_data_master_read;                                      // cpu1:d_read -> mm_interconnect_0:cpu1_data_master_read
	wire  [31:0] cpu1_data_master_readdata;                                  // mm_interconnect_0:cpu1_data_master_readdata -> cpu1:d_readdata
	wire         cpu1_data_master_debugaccess;                               // cpu1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu1_data_master_debugaccess
	wire   [3:0] cpu1_data_master_byteenable;                                // cpu1:d_byteenable -> mm_interconnect_0:cpu1_data_master_byteenable
	wire         cpu5_data_master_waitrequest;                               // mm_interconnect_0:cpu5_data_master_waitrequest -> cpu5:d_waitrequest
	wire  [31:0] cpu5_data_master_writedata;                                 // cpu5:d_writedata -> mm_interconnect_0:cpu5_data_master_writedata
	wire  [28:0] cpu5_data_master_address;                                   // cpu5:d_address -> mm_interconnect_0:cpu5_data_master_address
	wire         cpu5_data_master_write;                                     // cpu5:d_write -> mm_interconnect_0:cpu5_data_master_write
	wire         cpu5_data_master_read;                                      // cpu5:d_read -> mm_interconnect_0:cpu5_data_master_read
	wire  [31:0] cpu5_data_master_readdata;                                  // mm_interconnect_0:cpu5_data_master_readdata -> cpu5:d_readdata
	wire         cpu5_data_master_debugaccess;                               // cpu5:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu5_data_master_debugaccess
	wire   [3:0] cpu5_data_master_byteenable;                                // cpu5:d_byteenable -> mm_interconnect_0:cpu5_data_master_byteenable
	wire         cpu5_instruction_master_waitrequest;                        // mm_interconnect_0:cpu5_instruction_master_waitrequest -> cpu5:i_waitrequest
	wire  [17:0] cpu5_instruction_master_address;                            // cpu5:i_address -> mm_interconnect_0:cpu5_instruction_master_address
	wire         cpu5_instruction_master_read;                               // cpu5:i_read -> mm_interconnect_0:cpu5_instruction_master_read
	wire  [31:0] cpu5_instruction_master_readdata;                           // mm_interconnect_0:cpu5_instruction_master_readdata -> cpu5:i_readdata
	wire  [31:0] mm_interconnect_0_fifo1to6_in_csr_writedata;                // mm_interconnect_0:fifo1to6_in_csr_writedata -> fifo1to6:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo1to6_in_csr_address;                  // mm_interconnect_0:fifo1to6_in_csr_address -> fifo1to6:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo1to6_in_csr_write;                    // mm_interconnect_0:fifo1to6_in_csr_write -> fifo1to6:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo1to6_in_csr_read;                     // mm_interconnect_0:fifo1to6_in_csr_read -> fifo1to6:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to6_in_csr_readdata;                 // fifo1to6:wrclk_control_slave_readdata -> mm_interconnect_0:fifo1to6_in_csr_readdata
	wire  [31:0] mm_interconnect_0_fifo1to4_in_csr_writedata;                // mm_interconnect_0:fifo1to4_in_csr_writedata -> fifo1to4:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo1to4_in_csr_address;                  // mm_interconnect_0:fifo1to4_in_csr_address -> fifo1to4:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo1to4_in_csr_write;                    // mm_interconnect_0:fifo1to4_in_csr_write -> fifo1to4:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo1to4_in_csr_read;                     // mm_interconnect_0:fifo1to4_in_csr_read -> fifo1to4:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to4_in_csr_readdata;                 // fifo1to4:wrclk_control_slave_readdata -> mm_interconnect_0:fifo1to4_in_csr_readdata
	wire         cpu1_instruction_master_waitrequest;                        // mm_interconnect_0:cpu1_instruction_master_waitrequest -> cpu1:i_waitrequest
	wire  [28:0] cpu1_instruction_master_address;                            // cpu1:i_address -> mm_interconnect_0:cpu1_instruction_master_address
	wire         cpu1_instruction_master_read;                               // cpu1:i_read -> mm_interconnect_0:cpu1_instruction_master_read
	wire  [31:0] cpu1_instruction_master_readdata;                           // mm_interconnect_0:cpu1_instruction_master_readdata -> cpu1:i_readdata
	wire  [31:0] mm_interconnect_0_mem3_s1_writedata;                        // mm_interconnect_0:mem3_s1_writedata -> mem3:writedata
	wire  [14:0] mm_interconnect_0_mem3_s1_address;                          // mm_interconnect_0:mem3_s1_address -> mem3:address
	wire         mm_interconnect_0_mem3_s1_chipselect;                       // mm_interconnect_0:mem3_s1_chipselect -> mem3:chipselect
	wire         mm_interconnect_0_mem3_s1_clken;                            // mm_interconnect_0:mem3_s1_clken -> mem3:clken
	wire         mm_interconnect_0_mem3_s1_write;                            // mm_interconnect_0:mem3_s1_write -> mem3:write
	wire  [31:0] mm_interconnect_0_mem3_s1_readdata;                         // mem3:readdata -> mm_interconnect_0:mem3_s1_readdata
	wire   [3:0] mm_interconnect_0_mem3_s1_byteenable;                       // mm_interconnect_0:mem3_s1_byteenable -> mem3:byteenable
	wire  [31:0] mm_interconnect_0_mem6_s1_writedata;                        // mm_interconnect_0:mem6_s1_writedata -> mem6:writedata
	wire  [13:0] mm_interconnect_0_mem6_s1_address;                          // mm_interconnect_0:mem6_s1_address -> mem6:address
	wire         mm_interconnect_0_mem6_s1_chipselect;                       // mm_interconnect_0:mem6_s1_chipselect -> mem6:chipselect
	wire         mm_interconnect_0_mem6_s1_clken;                            // mm_interconnect_0:mem6_s1_clken -> mem6:clken
	wire         mm_interconnect_0_mem6_s1_write;                            // mm_interconnect_0:mem6_s1_write -> mem6:write
	wire  [31:0] mm_interconnect_0_mem6_s1_readdata;                         // mem6:readdata -> mm_interconnect_0:mem6_s1_readdata
	wire   [3:0] mm_interconnect_0_mem6_s1_byteenable;                       // mm_interconnect_0:mem6_s1_byteenable -> mem6:byteenable
	wire         mm_interconnect_0_fifo1to2a_in_waitrequest;                 // fifo1to2A:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo1to2A_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo1to2a_in_writedata;                   // mm_interconnect_0:fifo1to2A_in_writedata -> fifo1to2A:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo1to2a_in_write;                       // mm_interconnect_0:fifo1to2A_in_write -> fifo1to2A:avalonmm_write_slave_write
	wire         mm_interconnect_0_jtag_uart5_avalon_jtag_slave_waitrequest; // jtag_uart5:av_waitrequest -> mm_interconnect_0:jtag_uart5_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart5_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart5_avalon_jtag_slave_writedata -> jtag_uart5:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart5_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart5_avalon_jtag_slave_address -> jtag_uart5:av_address
	wire         mm_interconnect_0_jtag_uart5_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart5_avalon_jtag_slave_chipselect -> jtag_uart5:av_chipselect
	wire         mm_interconnect_0_jtag_uart5_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart5_avalon_jtag_slave_write -> jtag_uart5:av_write_n
	wire         mm_interconnect_0_jtag_uart5_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart5_avalon_jtag_slave_read -> jtag_uart5:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart5_avalon_jtag_slave_readdata;    // jtag_uart5:av_readdata -> mm_interconnect_0:jtag_uart5_avalon_jtag_slave_readdata
	wire         cpu6_instruction_master_waitrequest;                        // mm_interconnect_0:cpu6_instruction_master_waitrequest -> cpu6:i_waitrequest
	wire  [17:0] cpu6_instruction_master_address;                            // cpu6:i_address -> mm_interconnect_0:cpu6_instruction_master_address
	wire         cpu6_instruction_master_read;                               // cpu6:i_read -> mm_interconnect_0:cpu6_instruction_master_read
	wire  [31:0] cpu6_instruction_master_readdata;                           // mm_interconnect_0:cpu6_instruction_master_readdata -> cpu6:i_readdata
	wire         mm_interconnect_0_cpu6_jtag_debug_module_waitrequest;       // cpu6:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu6_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu6_jtag_debug_module_writedata;         // mm_interconnect_0:cpu6_jtag_debug_module_writedata -> cpu6:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu6_jtag_debug_module_address;           // mm_interconnect_0:cpu6_jtag_debug_module_address -> cpu6:jtag_debug_module_address
	wire         mm_interconnect_0_cpu6_jtag_debug_module_write;             // mm_interconnect_0:cpu6_jtag_debug_module_write -> cpu6:jtag_debug_module_write
	wire         mm_interconnect_0_cpu6_jtag_debug_module_read;              // mm_interconnect_0:cpu6_jtag_debug_module_read -> cpu6:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu6_jtag_debug_module_readdata;          // cpu6:jtag_debug_module_readdata -> mm_interconnect_0:cpu6_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu6_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu6_jtag_debug_module_debugaccess -> cpu6:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu6_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu6_jtag_debug_module_byteenable -> cpu6:jtag_debug_module_byteenable
	wire         cpu4_data_master_waitrequest;                               // mm_interconnect_0:cpu4_data_master_waitrequest -> cpu4:d_waitrequest
	wire  [31:0] cpu4_data_master_writedata;                                 // cpu4:d_writedata -> mm_interconnect_0:cpu4_data_master_writedata
	wire  [28:0] cpu4_data_master_address;                                   // cpu4:d_address -> mm_interconnect_0:cpu4_data_master_address
	wire         cpu4_data_master_write;                                     // cpu4:d_write -> mm_interconnect_0:cpu4_data_master_write
	wire         cpu4_data_master_read;                                      // cpu4:d_read -> mm_interconnect_0:cpu4_data_master_read
	wire  [31:0] cpu4_data_master_readdata;                                  // mm_interconnect_0:cpu4_data_master_readdata -> cpu4:d_readdata
	wire         cpu4_data_master_debugaccess;                               // cpu4:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu4_data_master_debugaccess
	wire   [3:0] cpu4_data_master_byteenable;                                // cpu4:d_byteenable -> mm_interconnect_0:cpu4_data_master_byteenable
	wire         mm_interconnect_0_cpu2_jtag_debug_module_waitrequest;       // cpu2:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu2_jtag_debug_module_writedata;         // mm_interconnect_0:cpu2_jtag_debug_module_writedata -> cpu2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu2_jtag_debug_module_address;           // mm_interconnect_0:cpu2_jtag_debug_module_address -> cpu2:jtag_debug_module_address
	wire         mm_interconnect_0_cpu2_jtag_debug_module_write;             // mm_interconnect_0:cpu2_jtag_debug_module_write -> cpu2:jtag_debug_module_write
	wire         mm_interconnect_0_cpu2_jtag_debug_module_read;              // mm_interconnect_0:cpu2_jtag_debug_module_read -> cpu2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu2_jtag_debug_module_readdata;          // cpu2:jtag_debug_module_readdata -> mm_interconnect_0:cpu2_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu2_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu2_jtag_debug_module_debugaccess -> cpu2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu2_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu2_jtag_debug_module_byteenable -> cpu2:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo1to6_in_waitrequest;                  // fifo1to6:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo1to6_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo1to6_in_writedata;                    // mm_interconnect_0:fifo1to6_in_writedata -> fifo1to6:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo1to6_in_write;                        // mm_interconnect_0:fifo1to6_in_write -> fifo1to6:avalonmm_write_slave_write
	wire         mm_interconnect_0_jtag_uart6_avalon_jtag_slave_waitrequest; // jtag_uart6:av_waitrequest -> mm_interconnect_0:jtag_uart6_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart6_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart6_avalon_jtag_slave_writedata -> jtag_uart6:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart6_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart6_avalon_jtag_slave_address -> jtag_uart6:av_address
	wire         mm_interconnect_0_jtag_uart6_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart6_avalon_jtag_slave_chipselect -> jtag_uart6:av_chipselect
	wire         mm_interconnect_0_jtag_uart6_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart6_avalon_jtag_slave_write -> jtag_uart6:av_write_n
	wire         mm_interconnect_0_jtag_uart6_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart6_avalon_jtag_slave_read -> jtag_uart6:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart6_avalon_jtag_slave_readdata;    // jtag_uart6:av_readdata -> mm_interconnect_0:jtag_uart6_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_fifo1to5_in_csr_writedata;                // mm_interconnect_0:fifo1to5_in_csr_writedata -> fifo1to5:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo1to5_in_csr_address;                  // mm_interconnect_0:fifo1to5_in_csr_address -> fifo1to5:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo1to5_in_csr_write;                    // mm_interconnect_0:fifo1to5_in_csr_write -> fifo1to5:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo1to5_in_csr_read;                     // mm_interconnect_0:fifo1to5_in_csr_read -> fifo1to5:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to5_in_csr_readdata;                 // fifo1to5:wrclk_control_slave_readdata -> mm_interconnect_0:fifo1to5_in_csr_readdata
	wire         mm_interconnect_0_jtag_uart3_avalon_jtag_slave_waitrequest; // jtag_uart3:av_waitrequest -> mm_interconnect_0:jtag_uart3_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart3_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart3_avalon_jtag_slave_writedata -> jtag_uart3:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart3_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart3_avalon_jtag_slave_address -> jtag_uart3:av_address
	wire         mm_interconnect_0_jtag_uart3_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart3_avalon_jtag_slave_chipselect -> jtag_uart3:av_chipselect
	wire         mm_interconnect_0_jtag_uart3_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart3_avalon_jtag_slave_write -> jtag_uart3:av_write_n
	wire         mm_interconnect_0_jtag_uart3_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart3_avalon_jtag_slave_read -> jtag_uart3:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart3_avalon_jtag_slave_readdata;    // jtag_uart3:av_readdata -> mm_interconnect_0:jtag_uart3_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_fifo4to5_in_csr_writedata;                // mm_interconnect_0:fifo4to5_in_csr_writedata -> fifo4to5:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo4to5_in_csr_address;                  // mm_interconnect_0:fifo4to5_in_csr_address -> fifo4to5:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo4to5_in_csr_write;                    // mm_interconnect_0:fifo4to5_in_csr_write -> fifo4to5:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo4to5_in_csr_read;                     // mm_interconnect_0:fifo4to5_in_csr_read -> fifo4to5:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo4to5_in_csr_readdata;                 // fifo4to5:wrclk_control_slave_readdata -> mm_interconnect_0:fifo4to5_in_csr_readdata
	wire         cpu3_data_master_waitrequest;                               // mm_interconnect_0:cpu3_data_master_waitrequest -> cpu3:d_waitrequest
	wire  [31:0] cpu3_data_master_writedata;                                 // cpu3:d_writedata -> mm_interconnect_0:cpu3_data_master_writedata
	wire  [28:0] cpu3_data_master_address;                                   // cpu3:d_address -> mm_interconnect_0:cpu3_data_master_address
	wire         cpu3_data_master_write;                                     // cpu3:d_write -> mm_interconnect_0:cpu3_data_master_write
	wire         cpu3_data_master_read;                                      // cpu3:d_read -> mm_interconnect_0:cpu3_data_master_read
	wire  [31:0] cpu3_data_master_readdata;                                  // mm_interconnect_0:cpu3_data_master_readdata -> cpu3:d_readdata
	wire         cpu3_data_master_debugaccess;                               // cpu3:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu3_data_master_debugaccess
	wire   [3:0] cpu3_data_master_byteenable;                                // cpu3:d_byteenable -> mm_interconnect_0:cpu3_data_master_byteenable
	wire         mm_interconnect_0_fifo1to4_out_waitrequest;                 // fifo1to4:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1to4_out_waitrequest
	wire         mm_interconnect_0_fifo1to4_out_read;                        // mm_interconnect_0:fifo1to4_out_read -> fifo1to4:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to4_out_readdata;                    // fifo1to4:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1to4_out_readdata
	wire         mm_interconnect_0_fifo1to2c_in_waitrequest;                 // fifo1to2C:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo1to2C_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo1to2c_in_writedata;                   // mm_interconnect_0:fifo1to2C_in_writedata -> fifo1to2C:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo1to2c_in_write;                       // mm_interconnect_0:fifo1to2C_in_write -> fifo1to2C:avalonmm_write_slave_write
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;              // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;             // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire  [31:0] mm_interconnect_0_mem4_s1_writedata;                        // mm_interconnect_0:mem4_s1_writedata -> mem4:writedata
	wire  [13:0] mm_interconnect_0_mem4_s1_address;                          // mm_interconnect_0:mem4_s1_address -> mem4:address
	wire         mm_interconnect_0_mem4_s1_chipselect;                       // mm_interconnect_0:mem4_s1_chipselect -> mem4:chipselect
	wire         mm_interconnect_0_mem4_s1_clken;                            // mm_interconnect_0:mem4_s1_clken -> mem4:clken
	wire         mm_interconnect_0_mem4_s1_write;                            // mm_interconnect_0:mem4_s1_write -> mem4:write
	wire  [31:0] mm_interconnect_0_mem4_s1_readdata;                         // mem4:readdata -> mm_interconnect_0:mem4_s1_readdata
	wire   [3:0] mm_interconnect_0_mem4_s1_byteenable;                       // mm_interconnect_0:mem4_s1_byteenable -> mem4:byteenable
	wire         cpu2_instruction_master_waitrequest;                        // mm_interconnect_0:cpu2_instruction_master_waitrequest -> cpu2:i_waitrequest
	wire  [18:0] cpu2_instruction_master_address;                            // cpu2:i_address -> mm_interconnect_0:cpu2_instruction_master_address
	wire         cpu2_instruction_master_read;                               // cpu2:i_read -> mm_interconnect_0:cpu2_instruction_master_read
	wire  [31:0] cpu2_instruction_master_readdata;                           // mm_interconnect_0:cpu2_instruction_master_readdata -> cpu2:i_readdata
	wire         mm_interconnect_0_cpu4_jtag_debug_module_waitrequest;       // cpu4:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu4_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu4_jtag_debug_module_writedata;         // mm_interconnect_0:cpu4_jtag_debug_module_writedata -> cpu4:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu4_jtag_debug_module_address;           // mm_interconnect_0:cpu4_jtag_debug_module_address -> cpu4:jtag_debug_module_address
	wire         mm_interconnect_0_cpu4_jtag_debug_module_write;             // mm_interconnect_0:cpu4_jtag_debug_module_write -> cpu4:jtag_debug_module_write
	wire         mm_interconnect_0_cpu4_jtag_debug_module_read;              // mm_interconnect_0:cpu4_jtag_debug_module_read -> cpu4:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu4_jtag_debug_module_readdata;          // cpu4:jtag_debug_module_readdata -> mm_interconnect_0:cpu4_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu4_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu4_jtag_debug_module_debugaccess -> cpu4:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu4_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu4_jtag_debug_module_byteenable -> cpu4:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo1to2a_out_waitrequest;                // fifo1to2A:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1to2A_out_waitrequest
	wire         mm_interconnect_0_fifo1to2a_out_read;                       // mm_interconnect_0:fifo1to2A_out_read -> fifo1to2A:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to2a_out_readdata;                   // fifo1to2A:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1to2A_out_readdata
	wire  [31:0] mm_interconnect_0_fifo5to6_in_csr_writedata;                // mm_interconnect_0:fifo5to6_in_csr_writedata -> fifo5to6:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo5to6_in_csr_address;                  // mm_interconnect_0:fifo5to6_in_csr_address -> fifo5to6:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo5to6_in_csr_write;                    // mm_interconnect_0:fifo5to6_in_csr_write -> fifo5to6:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo5to6_in_csr_read;                     // mm_interconnect_0:fifo5to6_in_csr_read -> fifo5to6:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo5to6_in_csr_readdata;                 // fifo5to6:wrclk_control_slave_readdata -> mm_interconnect_0:fifo5to6_in_csr_readdata
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest; // jtag_uart1:av_waitrequest -> mm_interconnect_0:jtag_uart1_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_writedata -> jtag_uart1:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_address -> jtag_uart1:av_address
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_chipselect -> jtag_uart1:av_chipselect
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_write -> jtag_uart1:av_write_n
	wire         mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart1_avalon_jtag_slave_read -> jtag_uart1:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata;    // jtag_uart1:av_readdata -> mm_interconnect_0:jtag_uart1_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_fifo3to4_in_csr_writedata;                // mm_interconnect_0:fifo3to4_in_csr_writedata -> fifo3to4:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo3to4_in_csr_address;                  // mm_interconnect_0:fifo3to4_in_csr_address -> fifo3to4:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo3to4_in_csr_write;                    // mm_interconnect_0:fifo3to4_in_csr_write -> fifo3to4:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo3to4_in_csr_read;                     // mm_interconnect_0:fifo3to4_in_csr_read -> fifo3to4:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo3to4_in_csr_readdata;                 // fifo3to4:wrclk_control_slave_readdata -> mm_interconnect_0:fifo3to4_in_csr_readdata
	wire  [15:0] mm_interconnect_0_timer1_s1_writedata;                      // mm_interconnect_0:timer1_s1_writedata -> timer1:writedata
	wire   [2:0] mm_interconnect_0_timer1_s1_address;                        // mm_interconnect_0:timer1_s1_address -> timer1:address
	wire         mm_interconnect_0_timer1_s1_chipselect;                     // mm_interconnect_0:timer1_s1_chipselect -> timer1:chipselect
	wire         mm_interconnect_0_timer1_s1_write;                          // mm_interconnect_0:timer1_s1_write -> timer1:write_n
	wire  [15:0] mm_interconnect_0_timer1_s1_readdata;                       // timer1:readdata -> mm_interconnect_0:timer1_s1_readdata
	wire         cpu3_instruction_master_waitrequest;                        // mm_interconnect_0:cpu3_instruction_master_waitrequest -> cpu3:i_waitrequest
	wire  [18:0] cpu3_instruction_master_address;                            // cpu3:i_address -> mm_interconnect_0:cpu3_instruction_master_address
	wire         cpu3_instruction_master_read;                               // cpu3:i_read -> mm_interconnect_0:cpu3_instruction_master_read
	wire  [31:0] cpu3_instruction_master_readdata;                           // mm_interconnect_0:cpu3_instruction_master_readdata -> cpu3:i_readdata
	wire  [31:0] mm_interconnect_0_fifo1to2b_in_csr_writedata;               // mm_interconnect_0:fifo1to2B_in_csr_writedata -> fifo1to2B:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo1to2b_in_csr_address;                 // mm_interconnect_0:fifo1to2B_in_csr_address -> fifo1to2B:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo1to2b_in_csr_write;                   // mm_interconnect_0:fifo1to2B_in_csr_write -> fifo1to2B:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo1to2b_in_csr_read;                    // mm_interconnect_0:fifo1to2B_in_csr_read -> fifo1to2B:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to2b_in_csr_readdata;                // fifo1to2B:wrclk_control_slave_readdata -> mm_interconnect_0:fifo1to2B_in_csr_readdata
	wire         mm_interconnect_0_cpu1_jtag_debug_module_waitrequest;       // cpu1:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu1_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu1_jtag_debug_module_writedata;         // mm_interconnect_0:cpu1_jtag_debug_module_writedata -> cpu1:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu1_jtag_debug_module_address;           // mm_interconnect_0:cpu1_jtag_debug_module_address -> cpu1:jtag_debug_module_address
	wire         mm_interconnect_0_cpu1_jtag_debug_module_write;             // mm_interconnect_0:cpu1_jtag_debug_module_write -> cpu1:jtag_debug_module_write
	wire         mm_interconnect_0_cpu1_jtag_debug_module_read;              // mm_interconnect_0:cpu1_jtag_debug_module_read -> cpu1:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu1_jtag_debug_module_readdata;          // cpu1:jtag_debug_module_readdata -> mm_interconnect_0:cpu1_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu1_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu1_jtag_debug_module_debugaccess -> cpu1:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu1_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu1_jtag_debug_module_byteenable -> cpu1:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo2to3_in_waitrequest;                  // fifo2to3:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo2to3_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo2to3_in_writedata;                    // mm_interconnect_0:fifo2to3_in_writedata -> fifo2to3:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo2to3_in_write;                        // mm_interconnect_0:fifo2to3_in_write -> fifo2to3:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_fifo2to3_in_csr_writedata;                // mm_interconnect_0:fifo2to3_in_csr_writedata -> fifo2to3:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo2to3_in_csr_address;                  // mm_interconnect_0:fifo2to3_in_csr_address -> fifo2to3:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo2to3_in_csr_write;                    // mm_interconnect_0:fifo2to3_in_csr_write -> fifo2to3:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo2to3_in_csr_read;                     // mm_interconnect_0:fifo2to3_in_csr_read -> fifo2to3:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo2to3_in_csr_readdata;                 // fifo2to3:wrclk_control_slave_readdata -> mm_interconnect_0:fifo2to3_in_csr_readdata
	wire  [15:0] mm_interconnect_0_timer5_s1_writedata;                      // mm_interconnect_0:timer5_s1_writedata -> timer5:writedata
	wire   [2:0] mm_interconnect_0_timer5_s1_address;                        // mm_interconnect_0:timer5_s1_address -> timer5:address
	wire         mm_interconnect_0_timer5_s1_chipselect;                     // mm_interconnect_0:timer5_s1_chipselect -> timer5:chipselect
	wire         mm_interconnect_0_timer5_s1_write;                          // mm_interconnect_0:timer5_s1_write -> timer5:write_n
	wire  [15:0] mm_interconnect_0_timer5_s1_readdata;                       // timer5:readdata -> mm_interconnect_0:timer5_s1_readdata
	wire         mm_interconnect_0_cpu3_jtag_debug_module_waitrequest;       // cpu3:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu3_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu3_jtag_debug_module_writedata;         // mm_interconnect_0:cpu3_jtag_debug_module_writedata -> cpu3:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu3_jtag_debug_module_address;           // mm_interconnect_0:cpu3_jtag_debug_module_address -> cpu3:jtag_debug_module_address
	wire         mm_interconnect_0_cpu3_jtag_debug_module_write;             // mm_interconnect_0:cpu3_jtag_debug_module_write -> cpu3:jtag_debug_module_write
	wire         mm_interconnect_0_cpu3_jtag_debug_module_read;              // mm_interconnect_0:cpu3_jtag_debug_module_read -> cpu3:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu3_jtag_debug_module_readdata;          // cpu3:jtag_debug_module_readdata -> mm_interconnect_0:cpu3_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu3_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu3_jtag_debug_module_debugaccess -> cpu3:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu3_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu3_jtag_debug_module_byteenable -> cpu3:jtag_debug_module_byteenable
	wire         mm_interconnect_0_fifo1to2b_in_waitrequest;                 // fifo1to2B:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo1to2B_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo1to2b_in_writedata;                   // mm_interconnect_0:fifo1to2B_in_writedata -> fifo1to2B:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo1to2b_in_write;                       // mm_interconnect_0:fifo1to2B_in_write -> fifo1to2B:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo5to6_in_waitrequest;                  // fifo5to6:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo5to6_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo5to6_in_writedata;                    // mm_interconnect_0:fifo5to6_in_writedata -> fifo5to6:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo5to6_in_write;                        // mm_interconnect_0:fifo5to6_in_write -> fifo5to6:avalonmm_write_slave_write
	wire         mm_interconnect_0_cpu5_jtag_debug_module_waitrequest;       // cpu5:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu5_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu5_jtag_debug_module_writedata;         // mm_interconnect_0:cpu5_jtag_debug_module_writedata -> cpu5:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu5_jtag_debug_module_address;           // mm_interconnect_0:cpu5_jtag_debug_module_address -> cpu5:jtag_debug_module_address
	wire         mm_interconnect_0_cpu5_jtag_debug_module_write;             // mm_interconnect_0:cpu5_jtag_debug_module_write -> cpu5:jtag_debug_module_write
	wire         mm_interconnect_0_cpu5_jtag_debug_module_read;              // mm_interconnect_0:cpu5_jtag_debug_module_read -> cpu5:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu5_jtag_debug_module_readdata;          // cpu5:jtag_debug_module_readdata -> mm_interconnect_0:cpu5_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu5_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu5_jtag_debug_module_debugaccess -> cpu5:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu5_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu5_jtag_debug_module_byteenable -> cpu5:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_fifo1to2c_in_csr_writedata;               // mm_interconnect_0:fifo1to2C_in_csr_writedata -> fifo1to2C:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo1to2c_in_csr_address;                 // mm_interconnect_0:fifo1to2C_in_csr_address -> fifo1to2C:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo1to2c_in_csr_write;                   // mm_interconnect_0:fifo1to2C_in_csr_write -> fifo1to2C:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo1to2c_in_csr_read;                    // mm_interconnect_0:fifo1to2C_in_csr_read -> fifo1to2C:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to2c_in_csr_readdata;                // fifo1to2C:wrclk_control_slave_readdata -> mm_interconnect_0:fifo1to2C_in_csr_readdata
	wire  [15:0] mm_interconnect_0_timer3_s1_writedata;                      // mm_interconnect_0:timer3_s1_writedata -> timer3:writedata
	wire   [2:0] mm_interconnect_0_timer3_s1_address;                        // mm_interconnect_0:timer3_s1_address -> timer3:address
	wire         mm_interconnect_0_timer3_s1_chipselect;                     // mm_interconnect_0:timer3_s1_chipselect -> timer3:chipselect
	wire         mm_interconnect_0_timer3_s1_write;                          // mm_interconnect_0:timer3_s1_write -> timer3:write_n
	wire  [15:0] mm_interconnect_0_timer3_s1_readdata;                       // timer3:readdata -> mm_interconnect_0:timer3_s1_readdata
	wire         mm_interconnect_0_fifo4to5_out_waitrequest;                 // fifo4to5:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo4to5_out_waitrequest
	wire         mm_interconnect_0_fifo4to5_out_read;                        // mm_interconnect_0:fifo4to5_out_read -> fifo4to5:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo4to5_out_readdata;                    // fifo4to5:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo4to5_out_readdata
	wire         mm_interconnect_0_fifo2to3_out_waitrequest;                 // fifo2to3:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo2to3_out_waitrequest
	wire         mm_interconnect_0_fifo2to3_out_read;                        // mm_interconnect_0:fifo2to3_out_read -> fifo2to3:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo2to3_out_readdata;                    // fifo2to3:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo2to3_out_readdata
	wire  [15:0] mm_interconnect_0_timer6_s1_writedata;                      // mm_interconnect_0:timer6_s1_writedata -> timer6:writedata
	wire   [2:0] mm_interconnect_0_timer6_s1_address;                        // mm_interconnect_0:timer6_s1_address -> timer6:address
	wire         mm_interconnect_0_timer6_s1_chipselect;                     // mm_interconnect_0:timer6_s1_chipselect -> timer6:chipselect
	wire         mm_interconnect_0_timer6_s1_write;                          // mm_interconnect_0:timer6_s1_write -> timer6:write_n
	wire  [15:0] mm_interconnect_0_timer6_s1_readdata;                       // timer6:readdata -> mm_interconnect_0:timer6_s1_readdata
	wire         mm_interconnect_0_fifo1to2b_out_waitrequest;                // fifo1to2B:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo1to2B_out_waitrequest
	wire         mm_interconnect_0_fifo1to2b_out_read;                       // mm_interconnect_0:fifo1to2B_out_read -> fifo1to2B:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo1to2b_out_readdata;                   // fifo1to2B:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo1to2B_out_readdata
	wire         mm_interconnect_0_jtag_uart2_avalon_jtag_slave_waitrequest; // jtag_uart2:av_waitrequest -> mm_interconnect_0:jtag_uart2_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart2_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart2_avalon_jtag_slave_writedata -> jtag_uart2:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart2_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart2_avalon_jtag_slave_address -> jtag_uart2:av_address
	wire         mm_interconnect_0_jtag_uart2_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart2_avalon_jtag_slave_chipselect -> jtag_uart2:av_chipselect
	wire         mm_interconnect_0_jtag_uart2_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart2_avalon_jtag_slave_write -> jtag_uart2:av_write_n
	wire         mm_interconnect_0_jtag_uart2_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart2_avalon_jtag_slave_read -> jtag_uart2:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart2_avalon_jtag_slave_readdata;    // jtag_uart2:av_readdata -> mm_interconnect_0:jtag_uart2_avalon_jtag_slave_readdata
	wire         cpu6_data_master_waitrequest;                               // mm_interconnect_0:cpu6_data_master_waitrequest -> cpu6:d_waitrequest
	wire  [31:0] cpu6_data_master_writedata;                                 // cpu6:d_writedata -> mm_interconnect_0:cpu6_data_master_writedata
	wire  [28:0] cpu6_data_master_address;                                   // cpu6:d_address -> mm_interconnect_0:cpu6_data_master_address
	wire         cpu6_data_master_write;                                     // cpu6:d_write -> mm_interconnect_0:cpu6_data_master_write
	wire         cpu6_data_master_read;                                      // cpu6:d_read -> mm_interconnect_0:cpu6_data_master_read
	wire  [31:0] cpu6_data_master_readdata;                                  // mm_interconnect_0:cpu6_data_master_readdata -> cpu6:d_readdata
	wire         cpu6_data_master_debugaccess;                               // cpu6:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu6_data_master_debugaccess
	wire   [3:0] cpu6_data_master_byteenable;                                // cpu6:d_byteenable -> mm_interconnect_0:cpu6_data_master_byteenable
	wire  [31:0] mm_interconnect_0_mem5_s1_writedata;                        // mm_interconnect_0:mem5_s1_writedata -> mem5:writedata
	wire  [13:0] mm_interconnect_0_mem5_s1_address;                          // mm_interconnect_0:mem5_s1_address -> mem5:address
	wire         mm_interconnect_0_mem5_s1_chipselect;                       // mm_interconnect_0:mem5_s1_chipselect -> mem5:chipselect
	wire         mm_interconnect_0_mem5_s1_clken;                            // mm_interconnect_0:mem5_s1_clken -> mem5:clken
	wire         mm_interconnect_0_mem5_s1_write;                            // mm_interconnect_0:mem5_s1_write -> mem5:write
	wire  [31:0] mm_interconnect_0_mem5_s1_readdata;                         // mem5:readdata -> mm_interconnect_0:mem5_s1_readdata
	wire   [3:0] mm_interconnect_0_mem5_s1_byteenable;                       // mm_interconnect_0:mem5_s1_byteenable -> mem5:byteenable
	wire         mm_interconnect_0_jtag_uart4_avalon_jtag_slave_waitrequest; // jtag_uart4:av_waitrequest -> mm_interconnect_0:jtag_uart4_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart4_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart4_avalon_jtag_slave_writedata -> jtag_uart4:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart4_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart4_avalon_jtag_slave_address -> jtag_uart4:av_address
	wire         mm_interconnect_0_jtag_uart4_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart4_avalon_jtag_slave_chipselect -> jtag_uart4:av_chipselect
	wire         mm_interconnect_0_jtag_uart4_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart4_avalon_jtag_slave_write -> jtag_uart4:av_write_n
	wire         mm_interconnect_0_jtag_uart4_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart4_avalon_jtag_slave_read -> jtag_uart4:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart4_avalon_jtag_slave_readdata;    // jtag_uart4:av_readdata -> mm_interconnect_0:jtag_uart4_avalon_jtag_slave_readdata
	wire         irq_mapper_receiver0_irq;                                   // timer1:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // jtag_uart1:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu1_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu1:d_irq
	wire         irq_mapper_001_receiver0_irq;                               // timer2:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                               // jtag_uart2:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] cpu2_d_irq_irq;                                             // irq_mapper_001:sender_irq -> cpu2:d_irq
	wire         irq_mapper_002_receiver0_irq;                               // timer3:irq -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                               // jtag_uart3:av_irq -> irq_mapper_002:receiver1_irq
	wire  [31:0] cpu3_d_irq_irq;                                             // irq_mapper_002:sender_irq -> cpu3:d_irq
	wire         irq_mapper_003_receiver0_irq;                               // timer4:irq -> irq_mapper_003:receiver0_irq
	wire         irq_mapper_003_receiver1_irq;                               // jtag_uart4:av_irq -> irq_mapper_003:receiver1_irq
	wire  [31:0] cpu4_d_irq_irq;                                             // irq_mapper_003:sender_irq -> cpu4:d_irq
	wire         irq_mapper_004_receiver0_irq;                               // timer5:irq -> irq_mapper_004:receiver0_irq
	wire         irq_mapper_004_receiver1_irq;                               // jtag_uart5:av_irq -> irq_mapper_004:receiver1_irq
	wire  [31:0] cpu5_d_irq_irq;                                             // irq_mapper_004:sender_irq -> cpu5:d_irq
	wire         irq_mapper_005_receiver0_irq;                               // timer6:irq -> irq_mapper_005:receiver0_irq
	wire         irq_mapper_005_receiver1_irq;                               // jtag_uart6:av_irq -> irq_mapper_005:receiver1_irq
	wire  [31:0] cpu6_d_irq_irq;                                             // irq_mapper_005:sender_irq -> cpu6:d_irq
	wire         irq_mapper_receiver2_irq;                                   // fifo1to2A:wrclk_control_slave_irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq]
	wire         irq_mapper_receiver3_irq;                                   // fifo1to2B:wrclk_control_slave_irq -> [irq_mapper:receiver3_irq, irq_mapper_001:receiver3_irq]
	wire         irq_mapper_receiver4_irq;                                   // fifo1to2C:wrclk_control_slave_irq -> [irq_mapper:receiver4_irq, irq_mapper_001:receiver4_irq]
	wire         irq_mapper_001_receiver5_irq;                               // fifo2to3:wrclk_control_slave_irq -> [irq_mapper_001:receiver5_irq, irq_mapper_002:receiver2_irq]
	wire         irq_mapper_002_receiver3_irq;                               // fifo3to4:wrclk_control_slave_irq -> [irq_mapper_002:receiver3_irq, irq_mapper_003:receiver2_irq]
	wire         irq_mapper_003_receiver3_irq;                               // fifo4to5:wrclk_control_slave_irq -> [irq_mapper_003:receiver3_irq, irq_mapper_004:receiver2_irq]
	wire         irq_mapper_004_receiver3_irq;                               // fifo5to6:wrclk_control_slave_irq -> [irq_mapper_004:receiver3_irq, irq_mapper_005:receiver2_irq]
	wire         irq_mapper_receiver5_irq;                                   // fifo1to4:wrclk_control_slave_irq -> [irq_mapper:receiver5_irq, irq_mapper_003:receiver4_irq]
	wire         irq_mapper_receiver6_irq;                                   // fifo1to5:wrclk_control_slave_irq -> [irq_mapper:receiver6_irq, irq_mapper_004:receiver4_irq]
	wire         irq_mapper_receiver7_irq;                                   // fifo1to6:wrclk_control_slave_irq -> [irq_mapper:receiver7_irq, irq_mapper_005:receiver3_irq]
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [cpu1:reset_n, irq_mapper:reset, jtag_uart1:rst_n, mm_interconnect_0:cpu1_reset_n_reset_bridge_in_reset_reset, pll:reset, rst_translator:in_reset, sdram_controller:reset_n, timer1:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [cpu1:reset_req, rst_translator:reset_req_in]
	wire         cpu1_jtag_debug_module_reset_reset;                         // cpu1:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_011:reset_in1, rst_controller_012:reset_in1, rst_controller_013:reset_in1, rst_controller_014:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [fifo1to2A:reset_n, fifo1to2B:reset_n, fifo1to2C:reset_n, mm_interconnect_0:fifo1to2A_reset_in_reset_bridge_in_reset_reset]
	wire         cpu2_jtag_debug_module_reset_reset;                         // cpu2:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in2, rst_controller_002:reset_in1, rst_controller_004:reset_in2, rst_controller_014:reset_in2]
	wire         rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [cpu2:reset_n, irq_mapper_001:reset, jtag_uart2:rst_n, mem2:reset, mm_interconnect_0:cpu2_reset_n_reset_bridge_in_reset_reset, rst_translator_001:in_reset, timer2:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                     // rst_controller_002:reset_req -> [cpu2:reset_req, mem2:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                         // rst_controller_003:reset_out -> [cpu3:reset_n, irq_mapper_002:reset, jtag_uart3:rst_n, mem3:reset, mm_interconnect_0:cpu3_reset_n_reset_bridge_in_reset_reset, rst_translator_002:in_reset, timer3:reset_n]
	wire         rst_controller_003_reset_out_reset_req;                     // rst_controller_003:reset_req -> [cpu3:reset_req, mem3:reset_req, rst_translator_002:reset_req_in]
	wire         cpu3_jtag_debug_module_reset_reset;                         // cpu3:jtag_debug_module_resetrequest -> [rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in0, rst_controller_014:reset_in3]
	wire         rst_controller_004_reset_out_reset;                         // rst_controller_004:reset_out -> [fifo2to3:reset_n, mm_interconnect_0:fifo2to3_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_005_reset_out_reset;                         // rst_controller_005:reset_out -> [fifo3to4:reset_n, mm_interconnect_0:fifo3to4_reset_in_reset_bridge_in_reset_reset]
	wire         cpu4_jtag_debug_module_reset_reset;                         // cpu4:jtag_debug_module_resetrequest -> [rst_controller_005:reset_in2, rst_controller_006:reset_in1, rst_controller_007:reset_in1, rst_controller_011:reset_in2, rst_controller_014:reset_in4]
	wire         rst_controller_006_reset_out_reset;                         // rst_controller_006:reset_out -> [cpu4:reset_n, irq_mapper_003:reset, jtag_uart4:rst_n, mem4:reset, mm_interconnect_0:cpu4_reset_n_reset_bridge_in_reset_reset, rst_translator_003:in_reset, timer4:reset_n]
	wire         rst_controller_006_reset_out_reset_req;                     // rst_controller_006:reset_req -> [cpu4:reset_req, mem4:reset_req, rst_translator_003:reset_req_in]
	wire         rst_controller_007_reset_out_reset;                         // rst_controller_007:reset_out -> [fifo4to5:reset_n, mm_interconnect_0:fifo4to5_reset_in_reset_bridge_in_reset_reset]
	wire         cpu5_jtag_debug_module_reset_reset;                         // cpu5:jtag_debug_module_resetrequest -> [rst_controller_007:reset_in2, rst_controller_008:reset_in1, rst_controller_009:reset_in0, rst_controller_012:reset_in2, rst_controller_014:reset_in5]
	wire         rst_controller_008_reset_out_reset;                         // rst_controller_008:reset_out -> [cpu5:reset_n, irq_mapper_004:reset, jtag_uart5:rst_n, mem5:reset, mm_interconnect_0:cpu5_reset_n_reset_bridge_in_reset_reset, rst_translator_004:in_reset, timer5:reset_n]
	wire         rst_controller_008_reset_out_reset_req;                     // rst_controller_008:reset_req -> [cpu5:reset_req, mem5:reset_req, rst_translator_004:reset_req_in]
	wire         rst_controller_009_reset_out_reset;                         // rst_controller_009:reset_out -> [fifo5to6:reset_n, mm_interconnect_0:fifo5to6_reset_in_reset_bridge_in_reset_reset]
	wire         cpu6_jtag_debug_module_reset_reset;                         // cpu6:jtag_debug_module_resetrequest -> [rst_controller_009:reset_in2, rst_controller_010:reset_in0, rst_controller_013:reset_in2, rst_controller_014:reset_in6]
	wire         rst_controller_010_reset_out_reset;                         // rst_controller_010:reset_out -> [cpu6:reset_n, irq_mapper_005:reset, jtag_uart6:rst_n, mem6:reset, mm_interconnect_0:cpu6_reset_n_reset_bridge_in_reset_reset, rst_translator_005:in_reset, timer6:reset_n]
	wire         rst_controller_010_reset_out_reset_req;                     // rst_controller_010:reset_req -> [cpu6:reset_req, mem6:reset_req, rst_translator_005:reset_req_in]
	wire         rst_controller_011_reset_out_reset;                         // rst_controller_011:reset_out -> [fifo1to4:reset_n, mm_interconnect_0:fifo1to4_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_012_reset_out_reset;                         // rst_controller_012:reset_out -> [fifo1to5:reset_n, mm_interconnect_0:fifo1to5_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_013_reset_out_reset;                         // rst_controller_013:reset_out -> [fifo1to6:reset_n, mm_interconnect_0:fifo1to6_reset_in_reset_bridge_in_reset_reset]
	wire         rst_controller_014_reset_out_reset;                         // rst_controller_014:reset_out -> [mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, sysid:reset_n]

	MSoC_cpu1 cpu1 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (cpu1_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu1_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu1_data_master_read),                                //                          .read
		.d_readdata                            (cpu1_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu1_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu1_data_master_write),                               //                          .write
		.d_writedata                           (cpu1_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu1_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu1_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu1_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu1_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu1_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu1_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu1_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu1_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu1_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu1_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu1_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu1_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu1_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu1_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu1_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	MSoC_timer1 timer1 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_0_timer1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                //   irq.irq
	);

	MSoC_jtag_uart1 jtag_uart1 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                            //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                    //               irq.irq
	);

	MSoC_fifo1to2A fifo1to2a (
		.wrclock                          (clk_clk),                                      //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),          // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo1to2a_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo1to2a_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo1to2a_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo1to2a_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo1to2a_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo1to2a_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo1to2a_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo1to2a_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo1to2a_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo1to2a_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo1to2a_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver2_irq)                      //   in_irq.irq
	);

	MSoC_fifo1to2A fifo1to2b (
		.wrclock                          (clk_clk),                                      //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),          // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo1to2b_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo1to2b_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo1to2b_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo1to2b_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo1to2b_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo1to2b_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo1to2b_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo1to2b_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo1to2b_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo1to2b_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo1to2b_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver3_irq)                      //   in_irq.irq
	);

	MSoC_fifo1to2A fifo1to2c (
		.wrclock                          (clk_clk),                                      //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),          // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo1to2c_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo1to2c_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo1to2c_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo1to2c_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo1to2c_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo1to2c_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo1to2c_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo1to2c_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo1to2c_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo1to2c_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo1to2c_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver4_irq)                      //   in_irq.irq
	);

	MSoC_cpu2 cpu2 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                  //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),               //                          .reset_req
		.d_address                             (cpu2_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu2_data_master_read),                                //                          .read
		.d_readdata                            (cpu2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu2_data_master_write),                               //                          .write
		.d_writedata                           (cpu2_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu2_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu2_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	MSoC_mem2 mem2 (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_mem2_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_mem2_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_mem2_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_mem2_s1_write),        //       .write
		.readdata   (mm_interconnect_0_mem2_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_mem2_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_mem2_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)  //       .reset_req
	);

	MSoC_timer1 timer2 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),    // reset.reset_n
		.address    (mm_interconnect_0_timer2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer2_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver0_irq)            //   irq.irq
	);

	MSoC_jtag_uart1 jtag_uart2 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart2_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart2_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                //               irq.irq
	);

	MSoC_cpu3 cpu3 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_003_reset_out_reset),                  //                   reset_n.reset_n
		.reset_req                             (rst_controller_003_reset_out_reset_req),               //                          .reset_req
		.d_address                             (cpu3_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu3_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu3_data_master_read),                                //                          .read
		.d_readdata                            (cpu3_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu3_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu3_data_master_write),                               //                          .write
		.d_writedata                           (cpu3_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu3_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu3_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu3_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu3_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu3_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu3_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu3_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu3_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu3_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu3_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu3_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu3_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu3_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu3_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu3_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	MSoC_mem3 mem3 (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_mem3_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_mem3_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_mem3_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_mem3_s1_write),        //       .write
		.readdata   (mm_interconnect_0_mem3_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_mem3_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_mem3_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req)  //       .reset_req
	);

	MSoC_timer1 timer3 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),    // reset.reset_n
		.address    (mm_interconnect_0_timer3_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer3_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer3_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer3_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer3_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver0_irq)            //   irq.irq
	);

	MSoC_jtag_uart1 jtag_uart3 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart3_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart3_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver1_irq)                                //               irq.irq
	);

	MSoC_fifo1to2A fifo2to3 (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_004_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo2to3_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo2to3_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo2to3_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo2to3_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo2to3_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo2to3_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo2to3_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo2to3_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo2to3_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo2to3_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo2to3_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_001_receiver5_irq)                 //   in_irq.irq
	);

	MSoC_fifo1to2A fifo3to4 (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_005_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo3to4_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo3to4_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo3to4_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo3to4_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo3to4_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo3to4_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo3to4_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo3to4_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo3to4_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo3to4_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo3to4_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_002_receiver3_irq)                 //   in_irq.irq
	);

	MSoC_cpu4 cpu4 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_006_reset_out_reset),                  //                   reset_n.reset_n
		.reset_req                             (rst_controller_006_reset_out_reset_req),               //                          .reset_req
		.d_address                             (cpu4_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu4_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu4_data_master_read),                                //                          .read
		.d_readdata                            (cpu4_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu4_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu4_data_master_write),                               //                          .write
		.d_writedata                           (cpu4_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu4_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu4_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu4_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu4_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu4_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu4_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu4_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu4_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu4_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu4_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu4_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu4_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu4_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu4_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu4_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	MSoC_mem4 mem4 (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_mem4_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_mem4_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_mem4_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_mem4_s1_write),        //       .write
		.readdata   (mm_interconnect_0_mem4_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_mem4_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_mem4_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_006_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_006_reset_out_reset_req)  //       .reset_req
	);

	MSoC_timer1 timer4 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_006_reset_out_reset),    // reset.reset_n
		.address    (mm_interconnect_0_timer4_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer4_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer4_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer4_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer4_s1_write),     //      .write_n
		.irq        (irq_mapper_003_receiver0_irq)            //   irq.irq
	);

	MSoC_jtag_uart1 jtag_uart4 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_006_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart4_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart4_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_003_receiver1_irq)                                //               irq.irq
	);

	MSoC_fifo1to2A fifo4to5 (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_007_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo4to5_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo4to5_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo4to5_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo4to5_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo4to5_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo4to5_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo4to5_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo4to5_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo4to5_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo4to5_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo4to5_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_003_receiver3_irq)                 //   in_irq.irq
	);

	MSoC_cpu5 cpu5 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_008_reset_out_reset),                  //                   reset_n.reset_n
		.reset_req                             (rst_controller_008_reset_out_reset_req),               //                          .reset_req
		.d_address                             (cpu5_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu5_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu5_data_master_read),                                //                          .read
		.d_readdata                            (cpu5_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu5_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu5_data_master_write),                               //                          .write
		.d_writedata                           (cpu5_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu5_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu5_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu5_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu5_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu5_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu5_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu5_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu5_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu5_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu5_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu5_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu5_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu5_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu5_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu5_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	MSoC_mem5 mem5 (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_mem5_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_mem5_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_mem5_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_mem5_s1_write),        //       .write
		.readdata   (mm_interconnect_0_mem5_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_mem5_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_mem5_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_008_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_008_reset_out_reset_req)  //       .reset_req
	);

	MSoC_timer1 timer5 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_008_reset_out_reset),    // reset.reset_n
		.address    (mm_interconnect_0_timer5_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer5_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer5_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer5_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer5_s1_write),     //      .write_n
		.irq        (irq_mapper_004_receiver0_irq)            //   irq.irq
	);

	MSoC_jtag_uart1 jtag_uart5 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_008_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart5_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart5_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_004_receiver1_irq)                                //               irq.irq
	);

	MSoC_fifo1to2A fifo5to6 (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_009_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo5to6_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo5to6_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo5to6_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo5to6_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo5to6_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo5to6_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo5to6_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo5to6_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo5to6_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo5to6_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo5to6_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_004_receiver3_irq)                 //   in_irq.irq
	);

	MSoC_cpu6 cpu6 (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_010_reset_out_reset),                  //                   reset_n.reset_n
		.reset_req                             (rst_controller_010_reset_out_reset_req),               //                          .reset_req
		.d_address                             (cpu6_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu6_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu6_data_master_read),                                //                          .read
		.d_readdata                            (cpu6_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu6_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu6_data_master_write),                               //                          .write
		.d_writedata                           (cpu6_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu6_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu6_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu6_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu6_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu6_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu6_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu6_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu6_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu6_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu6_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu6_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu6_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu6_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu6_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu6_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	MSoC_mem6 mem6 (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_mem6_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_mem6_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_mem6_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_mem6_s1_write),        //       .write
		.readdata   (mm_interconnect_0_mem6_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_mem6_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_mem6_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_010_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_010_reset_out_reset_req)  //       .reset_req
	);

	MSoC_timer1 timer6 (
		.clk        (clk_clk),                                //   clk.clk
		.reset_n    (~rst_controller_010_reset_out_reset),    // reset.reset_n
		.address    (mm_interconnect_0_timer6_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer6_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer6_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer6_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer6_s1_write),     //      .write_n
		.irq        (irq_mapper_005_receiver0_irq)            //   irq.irq
	);

	MSoC_jtag_uart1 jtag_uart6 (
		.clk            (clk_clk),                                                    //               clk.clk
		.rst_n          (~rst_controller_010_reset_out_reset),                        //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart6_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart6_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_005_receiver1_irq)                                //               irq.irq
	);

	MSoC_fifo1to2A fifo1to4 (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_011_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo1to4_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo1to4_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo1to4_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo1to4_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo1to4_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo1to4_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo1to4_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo1to4_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo1to4_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo1to4_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo1to4_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver5_irq)                     //   in_irq.irq
	);

	MSoC_fifo1to2A fifo1to5 (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_012_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo1to5_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo1to5_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo1to5_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo1to5_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo1to5_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo1to5_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo1to5_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo1to5_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo1to5_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo1to5_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo1to5_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver6_irq)                     //   in_irq.irq
	);

	MSoC_fifo1to2A fifo1to6 (
		.wrclock                          (clk_clk),                                     //   clk_in.clk
		.reset_n                          (~rst_controller_013_reset_out_reset),         // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo1to6_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo1to6_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo1to6_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo1to6_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo1to6_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo1to6_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo1to6_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo1to6_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo1to6_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo1to6_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo1to6_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver7_irq)                     //   in_irq.irq
	);

	MSoC_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_014_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	MSoC_sdram_controller sdram_controller (
		.clk            (clk_clk),                                             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	MSoC_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),            // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.areset    (),                                          //        areset_conduit.export
		.locked    (),                                          //        locked_conduit.export
		.phasedone ()                                           //     phasedone_conduit.export
	);

	MSoC_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                    (clk_clk),                                                    //                                  clk_clk.clk
		.cpu1_reset_n_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                             //       cpu1_reset_n_reset_bridge_in_reset.reset
		.cpu2_reset_n_reset_bridge_in_reset_reset       (rst_controller_002_reset_out_reset),                         //       cpu2_reset_n_reset_bridge_in_reset.reset
		.cpu3_reset_n_reset_bridge_in_reset_reset       (rst_controller_003_reset_out_reset),                         //       cpu3_reset_n_reset_bridge_in_reset.reset
		.cpu4_reset_n_reset_bridge_in_reset_reset       (rst_controller_006_reset_out_reset),                         //       cpu4_reset_n_reset_bridge_in_reset.reset
		.cpu5_reset_n_reset_bridge_in_reset_reset       (rst_controller_008_reset_out_reset),                         //       cpu5_reset_n_reset_bridge_in_reset.reset
		.cpu6_reset_n_reset_bridge_in_reset_reset       (rst_controller_010_reset_out_reset),                         //       cpu6_reset_n_reset_bridge_in_reset.reset
		.fifo1to2A_reset_in_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // fifo1to2A_reset_in_reset_bridge_in_reset.reset
		.fifo1to4_reset_in_reset_bridge_in_reset_reset  (rst_controller_011_reset_out_reset),                         //  fifo1to4_reset_in_reset_bridge_in_reset.reset
		.fifo1to5_reset_in_reset_bridge_in_reset_reset  (rst_controller_012_reset_out_reset),                         //  fifo1to5_reset_in_reset_bridge_in_reset.reset
		.fifo1to6_reset_in_reset_bridge_in_reset_reset  (rst_controller_013_reset_out_reset),                         //  fifo1to6_reset_in_reset_bridge_in_reset.reset
		.fifo2to3_reset_in_reset_bridge_in_reset_reset  (rst_controller_004_reset_out_reset),                         //  fifo2to3_reset_in_reset_bridge_in_reset.reset
		.fifo3to4_reset_in_reset_bridge_in_reset_reset  (rst_controller_005_reset_out_reset),                         //  fifo3to4_reset_in_reset_bridge_in_reset.reset
		.fifo4to5_reset_in_reset_bridge_in_reset_reset  (rst_controller_007_reset_out_reset),                         //  fifo4to5_reset_in_reset_bridge_in_reset.reset
		.fifo5to6_reset_in_reset_bridge_in_reset_reset  (rst_controller_009_reset_out_reset),                         //  fifo5to6_reset_in_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset        (rst_controller_014_reset_out_reset),                         //        sysid_reset_reset_bridge_in_reset.reset
		.cpu1_data_master_address                       (cpu1_data_master_address),                                   //                         cpu1_data_master.address
		.cpu1_data_master_waitrequest                   (cpu1_data_master_waitrequest),                               //                                         .waitrequest
		.cpu1_data_master_byteenable                    (cpu1_data_master_byteenable),                                //                                         .byteenable
		.cpu1_data_master_read                          (cpu1_data_master_read),                                      //                                         .read
		.cpu1_data_master_readdata                      (cpu1_data_master_readdata),                                  //                                         .readdata
		.cpu1_data_master_write                         (cpu1_data_master_write),                                     //                                         .write
		.cpu1_data_master_writedata                     (cpu1_data_master_writedata),                                 //                                         .writedata
		.cpu1_data_master_debugaccess                   (cpu1_data_master_debugaccess),                               //                                         .debugaccess
		.cpu1_instruction_master_address                (cpu1_instruction_master_address),                            //                  cpu1_instruction_master.address
		.cpu1_instruction_master_waitrequest            (cpu1_instruction_master_waitrequest),                        //                                         .waitrequest
		.cpu1_instruction_master_read                   (cpu1_instruction_master_read),                               //                                         .read
		.cpu1_instruction_master_readdata               (cpu1_instruction_master_readdata),                           //                                         .readdata
		.cpu2_data_master_address                       (cpu2_data_master_address),                                   //                         cpu2_data_master.address
		.cpu2_data_master_waitrequest                   (cpu2_data_master_waitrequest),                               //                                         .waitrequest
		.cpu2_data_master_byteenable                    (cpu2_data_master_byteenable),                                //                                         .byteenable
		.cpu2_data_master_read                          (cpu2_data_master_read),                                      //                                         .read
		.cpu2_data_master_readdata                      (cpu2_data_master_readdata),                                  //                                         .readdata
		.cpu2_data_master_write                         (cpu2_data_master_write),                                     //                                         .write
		.cpu2_data_master_writedata                     (cpu2_data_master_writedata),                                 //                                         .writedata
		.cpu2_data_master_debugaccess                   (cpu2_data_master_debugaccess),                               //                                         .debugaccess
		.cpu2_instruction_master_address                (cpu2_instruction_master_address),                            //                  cpu2_instruction_master.address
		.cpu2_instruction_master_waitrequest            (cpu2_instruction_master_waitrequest),                        //                                         .waitrequest
		.cpu2_instruction_master_read                   (cpu2_instruction_master_read),                               //                                         .read
		.cpu2_instruction_master_readdata               (cpu2_instruction_master_readdata),                           //                                         .readdata
		.cpu3_data_master_address                       (cpu3_data_master_address),                                   //                         cpu3_data_master.address
		.cpu3_data_master_waitrequest                   (cpu3_data_master_waitrequest),                               //                                         .waitrequest
		.cpu3_data_master_byteenable                    (cpu3_data_master_byteenable),                                //                                         .byteenable
		.cpu3_data_master_read                          (cpu3_data_master_read),                                      //                                         .read
		.cpu3_data_master_readdata                      (cpu3_data_master_readdata),                                  //                                         .readdata
		.cpu3_data_master_write                         (cpu3_data_master_write),                                     //                                         .write
		.cpu3_data_master_writedata                     (cpu3_data_master_writedata),                                 //                                         .writedata
		.cpu3_data_master_debugaccess                   (cpu3_data_master_debugaccess),                               //                                         .debugaccess
		.cpu3_instruction_master_address                (cpu3_instruction_master_address),                            //                  cpu3_instruction_master.address
		.cpu3_instruction_master_waitrequest            (cpu3_instruction_master_waitrequest),                        //                                         .waitrequest
		.cpu3_instruction_master_read                   (cpu3_instruction_master_read),                               //                                         .read
		.cpu3_instruction_master_readdata               (cpu3_instruction_master_readdata),                           //                                         .readdata
		.cpu4_data_master_address                       (cpu4_data_master_address),                                   //                         cpu4_data_master.address
		.cpu4_data_master_waitrequest                   (cpu4_data_master_waitrequest),                               //                                         .waitrequest
		.cpu4_data_master_byteenable                    (cpu4_data_master_byteenable),                                //                                         .byteenable
		.cpu4_data_master_read                          (cpu4_data_master_read),                                      //                                         .read
		.cpu4_data_master_readdata                      (cpu4_data_master_readdata),                                  //                                         .readdata
		.cpu4_data_master_write                         (cpu4_data_master_write),                                     //                                         .write
		.cpu4_data_master_writedata                     (cpu4_data_master_writedata),                                 //                                         .writedata
		.cpu4_data_master_debugaccess                   (cpu4_data_master_debugaccess),                               //                                         .debugaccess
		.cpu4_instruction_master_address                (cpu4_instruction_master_address),                            //                  cpu4_instruction_master.address
		.cpu4_instruction_master_waitrequest            (cpu4_instruction_master_waitrequest),                        //                                         .waitrequest
		.cpu4_instruction_master_read                   (cpu4_instruction_master_read),                               //                                         .read
		.cpu4_instruction_master_readdata               (cpu4_instruction_master_readdata),                           //                                         .readdata
		.cpu5_data_master_address                       (cpu5_data_master_address),                                   //                         cpu5_data_master.address
		.cpu5_data_master_waitrequest                   (cpu5_data_master_waitrequest),                               //                                         .waitrequest
		.cpu5_data_master_byteenable                    (cpu5_data_master_byteenable),                                //                                         .byteenable
		.cpu5_data_master_read                          (cpu5_data_master_read),                                      //                                         .read
		.cpu5_data_master_readdata                      (cpu5_data_master_readdata),                                  //                                         .readdata
		.cpu5_data_master_write                         (cpu5_data_master_write),                                     //                                         .write
		.cpu5_data_master_writedata                     (cpu5_data_master_writedata),                                 //                                         .writedata
		.cpu5_data_master_debugaccess                   (cpu5_data_master_debugaccess),                               //                                         .debugaccess
		.cpu5_instruction_master_address                (cpu5_instruction_master_address),                            //                  cpu5_instruction_master.address
		.cpu5_instruction_master_waitrequest            (cpu5_instruction_master_waitrequest),                        //                                         .waitrequest
		.cpu5_instruction_master_read                   (cpu5_instruction_master_read),                               //                                         .read
		.cpu5_instruction_master_readdata               (cpu5_instruction_master_readdata),                           //                                         .readdata
		.cpu6_data_master_address                       (cpu6_data_master_address),                                   //                         cpu6_data_master.address
		.cpu6_data_master_waitrequest                   (cpu6_data_master_waitrequest),                               //                                         .waitrequest
		.cpu6_data_master_byteenable                    (cpu6_data_master_byteenable),                                //                                         .byteenable
		.cpu6_data_master_read                          (cpu6_data_master_read),                                      //                                         .read
		.cpu6_data_master_readdata                      (cpu6_data_master_readdata),                                  //                                         .readdata
		.cpu6_data_master_write                         (cpu6_data_master_write),                                     //                                         .write
		.cpu6_data_master_writedata                     (cpu6_data_master_writedata),                                 //                                         .writedata
		.cpu6_data_master_debugaccess                   (cpu6_data_master_debugaccess),                               //                                         .debugaccess
		.cpu6_instruction_master_address                (cpu6_instruction_master_address),                            //                  cpu6_instruction_master.address
		.cpu6_instruction_master_waitrequest            (cpu6_instruction_master_waitrequest),                        //                                         .waitrequest
		.cpu6_instruction_master_read                   (cpu6_instruction_master_read),                               //                                         .read
		.cpu6_instruction_master_readdata               (cpu6_instruction_master_readdata),                           //                                         .readdata
		.cpu1_jtag_debug_module_address                 (mm_interconnect_0_cpu1_jtag_debug_module_address),           //                   cpu1_jtag_debug_module.address
		.cpu1_jtag_debug_module_write                   (mm_interconnect_0_cpu1_jtag_debug_module_write),             //                                         .write
		.cpu1_jtag_debug_module_read                    (mm_interconnect_0_cpu1_jtag_debug_module_read),              //                                         .read
		.cpu1_jtag_debug_module_readdata                (mm_interconnect_0_cpu1_jtag_debug_module_readdata),          //                                         .readdata
		.cpu1_jtag_debug_module_writedata               (mm_interconnect_0_cpu1_jtag_debug_module_writedata),         //                                         .writedata
		.cpu1_jtag_debug_module_byteenable              (mm_interconnect_0_cpu1_jtag_debug_module_byteenable),        //                                         .byteenable
		.cpu1_jtag_debug_module_waitrequest             (mm_interconnect_0_cpu1_jtag_debug_module_waitrequest),       //                                         .waitrequest
		.cpu1_jtag_debug_module_debugaccess             (mm_interconnect_0_cpu1_jtag_debug_module_debugaccess),       //                                         .debugaccess
		.cpu2_jtag_debug_module_address                 (mm_interconnect_0_cpu2_jtag_debug_module_address),           //                   cpu2_jtag_debug_module.address
		.cpu2_jtag_debug_module_write                   (mm_interconnect_0_cpu2_jtag_debug_module_write),             //                                         .write
		.cpu2_jtag_debug_module_read                    (mm_interconnect_0_cpu2_jtag_debug_module_read),              //                                         .read
		.cpu2_jtag_debug_module_readdata                (mm_interconnect_0_cpu2_jtag_debug_module_readdata),          //                                         .readdata
		.cpu2_jtag_debug_module_writedata               (mm_interconnect_0_cpu2_jtag_debug_module_writedata),         //                                         .writedata
		.cpu2_jtag_debug_module_byteenable              (mm_interconnect_0_cpu2_jtag_debug_module_byteenable),        //                                         .byteenable
		.cpu2_jtag_debug_module_waitrequest             (mm_interconnect_0_cpu2_jtag_debug_module_waitrequest),       //                                         .waitrequest
		.cpu2_jtag_debug_module_debugaccess             (mm_interconnect_0_cpu2_jtag_debug_module_debugaccess),       //                                         .debugaccess
		.cpu3_jtag_debug_module_address                 (mm_interconnect_0_cpu3_jtag_debug_module_address),           //                   cpu3_jtag_debug_module.address
		.cpu3_jtag_debug_module_write                   (mm_interconnect_0_cpu3_jtag_debug_module_write),             //                                         .write
		.cpu3_jtag_debug_module_read                    (mm_interconnect_0_cpu3_jtag_debug_module_read),              //                                         .read
		.cpu3_jtag_debug_module_readdata                (mm_interconnect_0_cpu3_jtag_debug_module_readdata),          //                                         .readdata
		.cpu3_jtag_debug_module_writedata               (mm_interconnect_0_cpu3_jtag_debug_module_writedata),         //                                         .writedata
		.cpu3_jtag_debug_module_byteenable              (mm_interconnect_0_cpu3_jtag_debug_module_byteenable),        //                                         .byteenable
		.cpu3_jtag_debug_module_waitrequest             (mm_interconnect_0_cpu3_jtag_debug_module_waitrequest),       //                                         .waitrequest
		.cpu3_jtag_debug_module_debugaccess             (mm_interconnect_0_cpu3_jtag_debug_module_debugaccess),       //                                         .debugaccess
		.cpu4_jtag_debug_module_address                 (mm_interconnect_0_cpu4_jtag_debug_module_address),           //                   cpu4_jtag_debug_module.address
		.cpu4_jtag_debug_module_write                   (mm_interconnect_0_cpu4_jtag_debug_module_write),             //                                         .write
		.cpu4_jtag_debug_module_read                    (mm_interconnect_0_cpu4_jtag_debug_module_read),              //                                         .read
		.cpu4_jtag_debug_module_readdata                (mm_interconnect_0_cpu4_jtag_debug_module_readdata),          //                                         .readdata
		.cpu4_jtag_debug_module_writedata               (mm_interconnect_0_cpu4_jtag_debug_module_writedata),         //                                         .writedata
		.cpu4_jtag_debug_module_byteenable              (mm_interconnect_0_cpu4_jtag_debug_module_byteenable),        //                                         .byteenable
		.cpu4_jtag_debug_module_waitrequest             (mm_interconnect_0_cpu4_jtag_debug_module_waitrequest),       //                                         .waitrequest
		.cpu4_jtag_debug_module_debugaccess             (mm_interconnect_0_cpu4_jtag_debug_module_debugaccess),       //                                         .debugaccess
		.cpu5_jtag_debug_module_address                 (mm_interconnect_0_cpu5_jtag_debug_module_address),           //                   cpu5_jtag_debug_module.address
		.cpu5_jtag_debug_module_write                   (mm_interconnect_0_cpu5_jtag_debug_module_write),             //                                         .write
		.cpu5_jtag_debug_module_read                    (mm_interconnect_0_cpu5_jtag_debug_module_read),              //                                         .read
		.cpu5_jtag_debug_module_readdata                (mm_interconnect_0_cpu5_jtag_debug_module_readdata),          //                                         .readdata
		.cpu5_jtag_debug_module_writedata               (mm_interconnect_0_cpu5_jtag_debug_module_writedata),         //                                         .writedata
		.cpu5_jtag_debug_module_byteenable              (mm_interconnect_0_cpu5_jtag_debug_module_byteenable),        //                                         .byteenable
		.cpu5_jtag_debug_module_waitrequest             (mm_interconnect_0_cpu5_jtag_debug_module_waitrequest),       //                                         .waitrequest
		.cpu5_jtag_debug_module_debugaccess             (mm_interconnect_0_cpu5_jtag_debug_module_debugaccess),       //                                         .debugaccess
		.cpu6_jtag_debug_module_address                 (mm_interconnect_0_cpu6_jtag_debug_module_address),           //                   cpu6_jtag_debug_module.address
		.cpu6_jtag_debug_module_write                   (mm_interconnect_0_cpu6_jtag_debug_module_write),             //                                         .write
		.cpu6_jtag_debug_module_read                    (mm_interconnect_0_cpu6_jtag_debug_module_read),              //                                         .read
		.cpu6_jtag_debug_module_readdata                (mm_interconnect_0_cpu6_jtag_debug_module_readdata),          //                                         .readdata
		.cpu6_jtag_debug_module_writedata               (mm_interconnect_0_cpu6_jtag_debug_module_writedata),         //                                         .writedata
		.cpu6_jtag_debug_module_byteenable              (mm_interconnect_0_cpu6_jtag_debug_module_byteenable),        //                                         .byteenable
		.cpu6_jtag_debug_module_waitrequest             (mm_interconnect_0_cpu6_jtag_debug_module_waitrequest),       //                                         .waitrequest
		.cpu6_jtag_debug_module_debugaccess             (mm_interconnect_0_cpu6_jtag_debug_module_debugaccess),       //                                         .debugaccess
		.fifo1to2A_in_write                             (mm_interconnect_0_fifo1to2a_in_write),                       //                             fifo1to2A_in.write
		.fifo1to2A_in_writedata                         (mm_interconnect_0_fifo1to2a_in_writedata),                   //                                         .writedata
		.fifo1to2A_in_waitrequest                       (mm_interconnect_0_fifo1to2a_in_waitrequest),                 //                                         .waitrequest
		.fifo1to2A_in_csr_address                       (mm_interconnect_0_fifo1to2a_in_csr_address),                 //                         fifo1to2A_in_csr.address
		.fifo1to2A_in_csr_write                         (mm_interconnect_0_fifo1to2a_in_csr_write),                   //                                         .write
		.fifo1to2A_in_csr_read                          (mm_interconnect_0_fifo1to2a_in_csr_read),                    //                                         .read
		.fifo1to2A_in_csr_readdata                      (mm_interconnect_0_fifo1to2a_in_csr_readdata),                //                                         .readdata
		.fifo1to2A_in_csr_writedata                     (mm_interconnect_0_fifo1to2a_in_csr_writedata),               //                                         .writedata
		.fifo1to2A_out_read                             (mm_interconnect_0_fifo1to2a_out_read),                       //                            fifo1to2A_out.read
		.fifo1to2A_out_readdata                         (mm_interconnect_0_fifo1to2a_out_readdata),                   //                                         .readdata
		.fifo1to2A_out_waitrequest                      (mm_interconnect_0_fifo1to2a_out_waitrequest),                //                                         .waitrequest
		.fifo1to2B_in_write                             (mm_interconnect_0_fifo1to2b_in_write),                       //                             fifo1to2B_in.write
		.fifo1to2B_in_writedata                         (mm_interconnect_0_fifo1to2b_in_writedata),                   //                                         .writedata
		.fifo1to2B_in_waitrequest                       (mm_interconnect_0_fifo1to2b_in_waitrequest),                 //                                         .waitrequest
		.fifo1to2B_in_csr_address                       (mm_interconnect_0_fifo1to2b_in_csr_address),                 //                         fifo1to2B_in_csr.address
		.fifo1to2B_in_csr_write                         (mm_interconnect_0_fifo1to2b_in_csr_write),                   //                                         .write
		.fifo1to2B_in_csr_read                          (mm_interconnect_0_fifo1to2b_in_csr_read),                    //                                         .read
		.fifo1to2B_in_csr_readdata                      (mm_interconnect_0_fifo1to2b_in_csr_readdata),                //                                         .readdata
		.fifo1to2B_in_csr_writedata                     (mm_interconnect_0_fifo1to2b_in_csr_writedata),               //                                         .writedata
		.fifo1to2B_out_read                             (mm_interconnect_0_fifo1to2b_out_read),                       //                            fifo1to2B_out.read
		.fifo1to2B_out_readdata                         (mm_interconnect_0_fifo1to2b_out_readdata),                   //                                         .readdata
		.fifo1to2B_out_waitrequest                      (mm_interconnect_0_fifo1to2b_out_waitrequest),                //                                         .waitrequest
		.fifo1to2C_in_write                             (mm_interconnect_0_fifo1to2c_in_write),                       //                             fifo1to2C_in.write
		.fifo1to2C_in_writedata                         (mm_interconnect_0_fifo1to2c_in_writedata),                   //                                         .writedata
		.fifo1to2C_in_waitrequest                       (mm_interconnect_0_fifo1to2c_in_waitrequest),                 //                                         .waitrequest
		.fifo1to2C_in_csr_address                       (mm_interconnect_0_fifo1to2c_in_csr_address),                 //                         fifo1to2C_in_csr.address
		.fifo1to2C_in_csr_write                         (mm_interconnect_0_fifo1to2c_in_csr_write),                   //                                         .write
		.fifo1to2C_in_csr_read                          (mm_interconnect_0_fifo1to2c_in_csr_read),                    //                                         .read
		.fifo1to2C_in_csr_readdata                      (mm_interconnect_0_fifo1to2c_in_csr_readdata),                //                                         .readdata
		.fifo1to2C_in_csr_writedata                     (mm_interconnect_0_fifo1to2c_in_csr_writedata),               //                                         .writedata
		.fifo1to2C_out_read                             (mm_interconnect_0_fifo1to2c_out_read),                       //                            fifo1to2C_out.read
		.fifo1to2C_out_readdata                         (mm_interconnect_0_fifo1to2c_out_readdata),                   //                                         .readdata
		.fifo1to2C_out_waitrequest                      (mm_interconnect_0_fifo1to2c_out_waitrequest),                //                                         .waitrequest
		.fifo1to4_in_write                              (mm_interconnect_0_fifo1to4_in_write),                        //                              fifo1to4_in.write
		.fifo1to4_in_writedata                          (mm_interconnect_0_fifo1to4_in_writedata),                    //                                         .writedata
		.fifo1to4_in_waitrequest                        (mm_interconnect_0_fifo1to4_in_waitrequest),                  //                                         .waitrequest
		.fifo1to4_in_csr_address                        (mm_interconnect_0_fifo1to4_in_csr_address),                  //                          fifo1to4_in_csr.address
		.fifo1to4_in_csr_write                          (mm_interconnect_0_fifo1to4_in_csr_write),                    //                                         .write
		.fifo1to4_in_csr_read                           (mm_interconnect_0_fifo1to4_in_csr_read),                     //                                         .read
		.fifo1to4_in_csr_readdata                       (mm_interconnect_0_fifo1to4_in_csr_readdata),                 //                                         .readdata
		.fifo1to4_in_csr_writedata                      (mm_interconnect_0_fifo1to4_in_csr_writedata),                //                                         .writedata
		.fifo1to4_out_read                              (mm_interconnect_0_fifo1to4_out_read),                        //                             fifo1to4_out.read
		.fifo1to4_out_readdata                          (mm_interconnect_0_fifo1to4_out_readdata),                    //                                         .readdata
		.fifo1to4_out_waitrequest                       (mm_interconnect_0_fifo1to4_out_waitrequest),                 //                                         .waitrequest
		.fifo1to5_in_write                              (mm_interconnect_0_fifo1to5_in_write),                        //                              fifo1to5_in.write
		.fifo1to5_in_writedata                          (mm_interconnect_0_fifo1to5_in_writedata),                    //                                         .writedata
		.fifo1to5_in_waitrequest                        (mm_interconnect_0_fifo1to5_in_waitrequest),                  //                                         .waitrequest
		.fifo1to5_in_csr_address                        (mm_interconnect_0_fifo1to5_in_csr_address),                  //                          fifo1to5_in_csr.address
		.fifo1to5_in_csr_write                          (mm_interconnect_0_fifo1to5_in_csr_write),                    //                                         .write
		.fifo1to5_in_csr_read                           (mm_interconnect_0_fifo1to5_in_csr_read),                     //                                         .read
		.fifo1to5_in_csr_readdata                       (mm_interconnect_0_fifo1to5_in_csr_readdata),                 //                                         .readdata
		.fifo1to5_in_csr_writedata                      (mm_interconnect_0_fifo1to5_in_csr_writedata),                //                                         .writedata
		.fifo1to5_out_read                              (mm_interconnect_0_fifo1to5_out_read),                        //                             fifo1to5_out.read
		.fifo1to5_out_readdata                          (mm_interconnect_0_fifo1to5_out_readdata),                    //                                         .readdata
		.fifo1to5_out_waitrequest                       (mm_interconnect_0_fifo1to5_out_waitrequest),                 //                                         .waitrequest
		.fifo1to6_in_write                              (mm_interconnect_0_fifo1to6_in_write),                        //                              fifo1to6_in.write
		.fifo1to6_in_writedata                          (mm_interconnect_0_fifo1to6_in_writedata),                    //                                         .writedata
		.fifo1to6_in_waitrequest                        (mm_interconnect_0_fifo1to6_in_waitrequest),                  //                                         .waitrequest
		.fifo1to6_in_csr_address                        (mm_interconnect_0_fifo1to6_in_csr_address),                  //                          fifo1to6_in_csr.address
		.fifo1to6_in_csr_write                          (mm_interconnect_0_fifo1to6_in_csr_write),                    //                                         .write
		.fifo1to6_in_csr_read                           (mm_interconnect_0_fifo1to6_in_csr_read),                     //                                         .read
		.fifo1to6_in_csr_readdata                       (mm_interconnect_0_fifo1to6_in_csr_readdata),                 //                                         .readdata
		.fifo1to6_in_csr_writedata                      (mm_interconnect_0_fifo1to6_in_csr_writedata),                //                                         .writedata
		.fifo1to6_out_read                              (mm_interconnect_0_fifo1to6_out_read),                        //                             fifo1to6_out.read
		.fifo1to6_out_readdata                          (mm_interconnect_0_fifo1to6_out_readdata),                    //                                         .readdata
		.fifo1to6_out_waitrequest                       (mm_interconnect_0_fifo1to6_out_waitrequest),                 //                                         .waitrequest
		.fifo2to3_in_write                              (mm_interconnect_0_fifo2to3_in_write),                        //                              fifo2to3_in.write
		.fifo2to3_in_writedata                          (mm_interconnect_0_fifo2to3_in_writedata),                    //                                         .writedata
		.fifo2to3_in_waitrequest                        (mm_interconnect_0_fifo2to3_in_waitrequest),                  //                                         .waitrequest
		.fifo2to3_in_csr_address                        (mm_interconnect_0_fifo2to3_in_csr_address),                  //                          fifo2to3_in_csr.address
		.fifo2to3_in_csr_write                          (mm_interconnect_0_fifo2to3_in_csr_write),                    //                                         .write
		.fifo2to3_in_csr_read                           (mm_interconnect_0_fifo2to3_in_csr_read),                     //                                         .read
		.fifo2to3_in_csr_readdata                       (mm_interconnect_0_fifo2to3_in_csr_readdata),                 //                                         .readdata
		.fifo2to3_in_csr_writedata                      (mm_interconnect_0_fifo2to3_in_csr_writedata),                //                                         .writedata
		.fifo2to3_out_read                              (mm_interconnect_0_fifo2to3_out_read),                        //                             fifo2to3_out.read
		.fifo2to3_out_readdata                          (mm_interconnect_0_fifo2to3_out_readdata),                    //                                         .readdata
		.fifo2to3_out_waitrequest                       (mm_interconnect_0_fifo2to3_out_waitrequest),                 //                                         .waitrequest
		.fifo3to4_in_write                              (mm_interconnect_0_fifo3to4_in_write),                        //                              fifo3to4_in.write
		.fifo3to4_in_writedata                          (mm_interconnect_0_fifo3to4_in_writedata),                    //                                         .writedata
		.fifo3to4_in_waitrequest                        (mm_interconnect_0_fifo3to4_in_waitrequest),                  //                                         .waitrequest
		.fifo3to4_in_csr_address                        (mm_interconnect_0_fifo3to4_in_csr_address),                  //                          fifo3to4_in_csr.address
		.fifo3to4_in_csr_write                          (mm_interconnect_0_fifo3to4_in_csr_write),                    //                                         .write
		.fifo3to4_in_csr_read                           (mm_interconnect_0_fifo3to4_in_csr_read),                     //                                         .read
		.fifo3to4_in_csr_readdata                       (mm_interconnect_0_fifo3to4_in_csr_readdata),                 //                                         .readdata
		.fifo3to4_in_csr_writedata                      (mm_interconnect_0_fifo3to4_in_csr_writedata),                //                                         .writedata
		.fifo3to4_out_read                              (mm_interconnect_0_fifo3to4_out_read),                        //                             fifo3to4_out.read
		.fifo3to4_out_readdata                          (mm_interconnect_0_fifo3to4_out_readdata),                    //                                         .readdata
		.fifo3to4_out_waitrequest                       (mm_interconnect_0_fifo3to4_out_waitrequest),                 //                                         .waitrequest
		.fifo4to5_in_write                              (mm_interconnect_0_fifo4to5_in_write),                        //                              fifo4to5_in.write
		.fifo4to5_in_writedata                          (mm_interconnect_0_fifo4to5_in_writedata),                    //                                         .writedata
		.fifo4to5_in_waitrequest                        (mm_interconnect_0_fifo4to5_in_waitrequest),                  //                                         .waitrequest
		.fifo4to5_in_csr_address                        (mm_interconnect_0_fifo4to5_in_csr_address),                  //                          fifo4to5_in_csr.address
		.fifo4to5_in_csr_write                          (mm_interconnect_0_fifo4to5_in_csr_write),                    //                                         .write
		.fifo4to5_in_csr_read                           (mm_interconnect_0_fifo4to5_in_csr_read),                     //                                         .read
		.fifo4to5_in_csr_readdata                       (mm_interconnect_0_fifo4to5_in_csr_readdata),                 //                                         .readdata
		.fifo4to5_in_csr_writedata                      (mm_interconnect_0_fifo4to5_in_csr_writedata),                //                                         .writedata
		.fifo4to5_out_read                              (mm_interconnect_0_fifo4to5_out_read),                        //                             fifo4to5_out.read
		.fifo4to5_out_readdata                          (mm_interconnect_0_fifo4to5_out_readdata),                    //                                         .readdata
		.fifo4to5_out_waitrequest                       (mm_interconnect_0_fifo4to5_out_waitrequest),                 //                                         .waitrequest
		.fifo5to6_in_write                              (mm_interconnect_0_fifo5to6_in_write),                        //                              fifo5to6_in.write
		.fifo5to6_in_writedata                          (mm_interconnect_0_fifo5to6_in_writedata),                    //                                         .writedata
		.fifo5to6_in_waitrequest                        (mm_interconnect_0_fifo5to6_in_waitrequest),                  //                                         .waitrequest
		.fifo5to6_in_csr_address                        (mm_interconnect_0_fifo5to6_in_csr_address),                  //                          fifo5to6_in_csr.address
		.fifo5to6_in_csr_write                          (mm_interconnect_0_fifo5to6_in_csr_write),                    //                                         .write
		.fifo5to6_in_csr_read                           (mm_interconnect_0_fifo5to6_in_csr_read),                     //                                         .read
		.fifo5to6_in_csr_readdata                       (mm_interconnect_0_fifo5to6_in_csr_readdata),                 //                                         .readdata
		.fifo5to6_in_csr_writedata                      (mm_interconnect_0_fifo5to6_in_csr_writedata),                //                                         .writedata
		.fifo5to6_out_read                              (mm_interconnect_0_fifo5to6_out_read),                        //                             fifo5to6_out.read
		.fifo5to6_out_readdata                          (mm_interconnect_0_fifo5to6_out_readdata),                    //                                         .readdata
		.fifo5to6_out_waitrequest                       (mm_interconnect_0_fifo5to6_out_waitrequest),                 //                                         .waitrequest
		.jtag_uart1_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_address),     //             jtag_uart1_avalon_jtag_slave.address
		.jtag_uart1_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart1_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart1_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart1_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart1_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart1_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart1_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.jtag_uart2_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_address),     //             jtag_uart2_avalon_jtag_slave.address
		.jtag_uart2_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart2_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart2_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart2_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart2_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart2_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart2_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.jtag_uart3_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_address),     //             jtag_uart3_avalon_jtag_slave.address
		.jtag_uart3_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart3_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart3_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart3_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart3_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart3_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart3_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.jtag_uart4_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_address),     //             jtag_uart4_avalon_jtag_slave.address
		.jtag_uart4_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart4_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart4_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart4_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart4_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart4_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart4_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.jtag_uart5_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_address),     //             jtag_uart5_avalon_jtag_slave.address
		.jtag_uart5_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart5_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart5_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart5_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart5_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart5_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart5_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.jtag_uart6_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_address),     //             jtag_uart6_avalon_jtag_slave.address
		.jtag_uart6_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart6_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart6_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart6_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart6_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart6_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart6_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.mem2_s1_address                                (mm_interconnect_0_mem2_s1_address),                          //                                  mem2_s1.address
		.mem2_s1_write                                  (mm_interconnect_0_mem2_s1_write),                            //                                         .write
		.mem2_s1_readdata                               (mm_interconnect_0_mem2_s1_readdata),                         //                                         .readdata
		.mem2_s1_writedata                              (mm_interconnect_0_mem2_s1_writedata),                        //                                         .writedata
		.mem2_s1_byteenable                             (mm_interconnect_0_mem2_s1_byteenable),                       //                                         .byteenable
		.mem2_s1_chipselect                             (mm_interconnect_0_mem2_s1_chipselect),                       //                                         .chipselect
		.mem2_s1_clken                                  (mm_interconnect_0_mem2_s1_clken),                            //                                         .clken
		.mem3_s1_address                                (mm_interconnect_0_mem3_s1_address),                          //                                  mem3_s1.address
		.mem3_s1_write                                  (mm_interconnect_0_mem3_s1_write),                            //                                         .write
		.mem3_s1_readdata                               (mm_interconnect_0_mem3_s1_readdata),                         //                                         .readdata
		.mem3_s1_writedata                              (mm_interconnect_0_mem3_s1_writedata),                        //                                         .writedata
		.mem3_s1_byteenable                             (mm_interconnect_0_mem3_s1_byteenable),                       //                                         .byteenable
		.mem3_s1_chipselect                             (mm_interconnect_0_mem3_s1_chipselect),                       //                                         .chipselect
		.mem3_s1_clken                                  (mm_interconnect_0_mem3_s1_clken),                            //                                         .clken
		.mem4_s1_address                                (mm_interconnect_0_mem4_s1_address),                          //                                  mem4_s1.address
		.mem4_s1_write                                  (mm_interconnect_0_mem4_s1_write),                            //                                         .write
		.mem4_s1_readdata                               (mm_interconnect_0_mem4_s1_readdata),                         //                                         .readdata
		.mem4_s1_writedata                              (mm_interconnect_0_mem4_s1_writedata),                        //                                         .writedata
		.mem4_s1_byteenable                             (mm_interconnect_0_mem4_s1_byteenable),                       //                                         .byteenable
		.mem4_s1_chipselect                             (mm_interconnect_0_mem4_s1_chipselect),                       //                                         .chipselect
		.mem4_s1_clken                                  (mm_interconnect_0_mem4_s1_clken),                            //                                         .clken
		.mem5_s1_address                                (mm_interconnect_0_mem5_s1_address),                          //                                  mem5_s1.address
		.mem5_s1_write                                  (mm_interconnect_0_mem5_s1_write),                            //                                         .write
		.mem5_s1_readdata                               (mm_interconnect_0_mem5_s1_readdata),                         //                                         .readdata
		.mem5_s1_writedata                              (mm_interconnect_0_mem5_s1_writedata),                        //                                         .writedata
		.mem5_s1_byteenable                             (mm_interconnect_0_mem5_s1_byteenable),                       //                                         .byteenable
		.mem5_s1_chipselect                             (mm_interconnect_0_mem5_s1_chipselect),                       //                                         .chipselect
		.mem5_s1_clken                                  (mm_interconnect_0_mem5_s1_clken),                            //                                         .clken
		.mem6_s1_address                                (mm_interconnect_0_mem6_s1_address),                          //                                  mem6_s1.address
		.mem6_s1_write                                  (mm_interconnect_0_mem6_s1_write),                            //                                         .write
		.mem6_s1_readdata                               (mm_interconnect_0_mem6_s1_readdata),                         //                                         .readdata
		.mem6_s1_writedata                              (mm_interconnect_0_mem6_s1_writedata),                        //                                         .writedata
		.mem6_s1_byteenable                             (mm_interconnect_0_mem6_s1_byteenable),                       //                                         .byteenable
		.mem6_s1_chipselect                             (mm_interconnect_0_mem6_s1_chipselect),                       //                                         .chipselect
		.mem6_s1_clken                                  (mm_interconnect_0_mem6_s1_clken),                            //                                         .clken
		.pll_pll_slave_address                          (mm_interconnect_0_pll_pll_slave_address),                    //                            pll_pll_slave.address
		.pll_pll_slave_write                            (mm_interconnect_0_pll_pll_slave_write),                      //                                         .write
		.pll_pll_slave_read                             (mm_interconnect_0_pll_pll_slave_read),                       //                                         .read
		.pll_pll_slave_readdata                         (mm_interconnect_0_pll_pll_slave_readdata),                   //                                         .readdata
		.pll_pll_slave_writedata                        (mm_interconnect_0_pll_pll_slave_writedata),                  //                                         .writedata
		.sdram_controller_s1_address                    (mm_interconnect_0_sdram_controller_s1_address),              //                      sdram_controller_s1.address
		.sdram_controller_s1_write                      (mm_interconnect_0_sdram_controller_s1_write),                //                                         .write
		.sdram_controller_s1_read                       (mm_interconnect_0_sdram_controller_s1_read),                 //                                         .read
		.sdram_controller_s1_readdata                   (mm_interconnect_0_sdram_controller_s1_readdata),             //                                         .readdata
		.sdram_controller_s1_writedata                  (mm_interconnect_0_sdram_controller_s1_writedata),            //                                         .writedata
		.sdram_controller_s1_byteenable                 (mm_interconnect_0_sdram_controller_s1_byteenable),           //                                         .byteenable
		.sdram_controller_s1_readdatavalid              (mm_interconnect_0_sdram_controller_s1_readdatavalid),        //                                         .readdatavalid
		.sdram_controller_s1_waitrequest                (mm_interconnect_0_sdram_controller_s1_waitrequest),          //                                         .waitrequest
		.sdram_controller_s1_chipselect                 (mm_interconnect_0_sdram_controller_s1_chipselect),           //                                         .chipselect
		.sysid_control_slave_address                    (mm_interconnect_0_sysid_control_slave_address),              //                      sysid_control_slave.address
		.sysid_control_slave_readdata                   (mm_interconnect_0_sysid_control_slave_readdata),             //                                         .readdata
		.timer1_s1_address                              (mm_interconnect_0_timer1_s1_address),                        //                                timer1_s1.address
		.timer1_s1_write                                (mm_interconnect_0_timer1_s1_write),                          //                                         .write
		.timer1_s1_readdata                             (mm_interconnect_0_timer1_s1_readdata),                       //                                         .readdata
		.timer1_s1_writedata                            (mm_interconnect_0_timer1_s1_writedata),                      //                                         .writedata
		.timer1_s1_chipselect                           (mm_interconnect_0_timer1_s1_chipselect),                     //                                         .chipselect
		.timer2_s1_address                              (mm_interconnect_0_timer2_s1_address),                        //                                timer2_s1.address
		.timer2_s1_write                                (mm_interconnect_0_timer2_s1_write),                          //                                         .write
		.timer2_s1_readdata                             (mm_interconnect_0_timer2_s1_readdata),                       //                                         .readdata
		.timer2_s1_writedata                            (mm_interconnect_0_timer2_s1_writedata),                      //                                         .writedata
		.timer2_s1_chipselect                           (mm_interconnect_0_timer2_s1_chipselect),                     //                                         .chipselect
		.timer3_s1_address                              (mm_interconnect_0_timer3_s1_address),                        //                                timer3_s1.address
		.timer3_s1_write                                (mm_interconnect_0_timer3_s1_write),                          //                                         .write
		.timer3_s1_readdata                             (mm_interconnect_0_timer3_s1_readdata),                       //                                         .readdata
		.timer3_s1_writedata                            (mm_interconnect_0_timer3_s1_writedata),                      //                                         .writedata
		.timer3_s1_chipselect                           (mm_interconnect_0_timer3_s1_chipselect),                     //                                         .chipselect
		.timer4_s1_address                              (mm_interconnect_0_timer4_s1_address),                        //                                timer4_s1.address
		.timer4_s1_write                                (mm_interconnect_0_timer4_s1_write),                          //                                         .write
		.timer4_s1_readdata                             (mm_interconnect_0_timer4_s1_readdata),                       //                                         .readdata
		.timer4_s1_writedata                            (mm_interconnect_0_timer4_s1_writedata),                      //                                         .writedata
		.timer4_s1_chipselect                           (mm_interconnect_0_timer4_s1_chipselect),                     //                                         .chipselect
		.timer5_s1_address                              (mm_interconnect_0_timer5_s1_address),                        //                                timer5_s1.address
		.timer5_s1_write                                (mm_interconnect_0_timer5_s1_write),                          //                                         .write
		.timer5_s1_readdata                             (mm_interconnect_0_timer5_s1_readdata),                       //                                         .readdata
		.timer5_s1_writedata                            (mm_interconnect_0_timer5_s1_writedata),                      //                                         .writedata
		.timer5_s1_chipselect                           (mm_interconnect_0_timer5_s1_chipselect),                     //                                         .chipselect
		.timer6_s1_address                              (mm_interconnect_0_timer6_s1_address),                        //                                timer6_s1.address
		.timer6_s1_write                                (mm_interconnect_0_timer6_s1_write),                          //                                         .write
		.timer6_s1_readdata                             (mm_interconnect_0_timer6_s1_readdata),                       //                                         .readdata
		.timer6_s1_writedata                            (mm_interconnect_0_timer6_s1_writedata),                      //                                         .writedata
		.timer6_s1_chipselect                           (mm_interconnect_0_timer6_s1_chipselect)                      //                                         .chipselect
	);

	MSoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.sender_irq    (cpu1_d_irq_irq)                  //    sender.irq
	);

	MSoC_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_001_receiver5_irq),       // receiver5.irq
		.sender_irq    (cpu2_d_irq_irq)                      //    sender.irq
	);

	MSoC_irq_mapper_002 irq_mapper_002 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_001_receiver5_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_002_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu3_d_irq_irq)                      //    sender.irq
	);

	MSoC_irq_mapper_003 irq_mapper_003 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_006_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_003_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_003_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_002_receiver3_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_003_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver5_irq),           // receiver4.irq
		.sender_irq    (cpu4_d_irq_irq)                      //    sender.irq
	);

	MSoC_irq_mapper_003 irq_mapper_004 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_008_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_004_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_004_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_003_receiver3_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_004_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver6_irq),           // receiver4.irq
		.sender_irq    (cpu5_d_irq_irq)                      //    sender.irq
	);

	MSoC_irq_mapper_002 irq_mapper_005 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_010_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_005_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_005_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_004_receiver3_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver7_irq),           // receiver3.irq
		.sender_irq    (cpu6_d_irq_irq)                      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu2_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu2_jtag_debug_module_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu3_jtag_debug_module_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu3_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu2_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (cpu3_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (cpu4_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu4_jtag_debug_module_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_006_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu4_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu5_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu5_jtag_debug_module_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_008_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_009 (
		.reset_in0      (cpu5_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (cpu6_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_009_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_010 (
		.reset_in0      (cpu6_jtag_debug_module_reset_reset),     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_010_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_010_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_011 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu4_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_011_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_012 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu5_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_012_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_013 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu6_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_013_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (7),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_014 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu2_jtag_debug_module_reset_reset), // reset_in2.reset
		.reset_in3      (cpu3_jtag_debug_module_reset_reset), // reset_in3.reset
		.reset_in4      (cpu4_jtag_debug_module_reset_reset), // reset_in4.reset
		.reset_in5      (cpu5_jtag_debug_module_reset_reset), // reset_in5.reset
		.reset_in6      (cpu6_jtag_debug_module_reset_reset), // reset_in6.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_014_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
